/******************************************************************************
*
*  Authors:   Chengyi Zhang
*     Date:   2023/4/20
*   Method:   
*  Version:   
*  Content:  
* 
******************************************************************************/

module img_buffer (
    input   [   4: 0]                   i_addr                     ,
    output  [   7: 0]                   o_data [  2: 0]  [ 27: 0]
);

logic [7:0] rom [27:0][27:0];

generate
    for (genvar i = 0; i < 3; i++) begin
        for (genvar j = 0; j < 28; j++) begin
            assign o_data[i][j] = rom[i_addr + i][j];
        end
    end
endgenerate

assign rom[0][0] = 0;
assign rom[0][1] = 0;
assign rom[0][2] = 0;
assign rom[0][3] = 0;
assign rom[0][4] = 0;
assign rom[0][5] = 0;
assign rom[0][6] = 0;
assign rom[0][7] = 0;
assign rom[0][8] = 0;
assign rom[0][9] = 0;
assign rom[0][10] = 0;
assign rom[0][11] = 0;
assign rom[0][12] = 0;
assign rom[0][13] = 0;
assign rom[0][14] = 0;
assign rom[0][15] = 0;
assign rom[0][16] = 0;
assign rom[0][17] = 0;
assign rom[0][18] = 0;
assign rom[0][19] = 0;
assign rom[0][20] = 0;
assign rom[0][21] = 0;
assign rom[0][22] = 0;
assign rom[0][23] = 0;
assign rom[0][24] = 0;
assign rom[0][25] = 0;
assign rom[0][26] = 0;
assign rom[0][27] = 0;
assign rom[1][0] = 0;
assign rom[1][1] = 0;
assign rom[1][2] = 0;
assign rom[1][3] = 0;
assign rom[1][4] = 0;
assign rom[1][5] = 0;
assign rom[1][6] = 0;
assign rom[1][7] = 0;
assign rom[1][8] = 0;
assign rom[1][9] = 0;
assign rom[1][10] = 0;
assign rom[1][11] = 0;
assign rom[1][12] = 0;
assign rom[1][13] = 0;
assign rom[1][14] = 0;
assign rom[1][15] = 0;
assign rom[1][16] = 0;
assign rom[1][17] = 0;
assign rom[1][18] = 0;
assign rom[1][19] = 0;
assign rom[1][20] = 0;
assign rom[1][21] = 0;
assign rom[1][22] = 0;
assign rom[1][23] = 0;
assign rom[1][24] = 0;
assign rom[1][25] = 0;
assign rom[1][26] = 0;
assign rom[1][27] = 0;
assign rom[2][0] = 0;
assign rom[2][1] = 0;
assign rom[2][2] = 0;
assign rom[2][3] = 0;
assign rom[2][4] = 0;
assign rom[2][5] = 0;
assign rom[2][6] = 0;
assign rom[2][7] = 0;
assign rom[2][8] = 0;
assign rom[2][9] = 0;
assign rom[2][10] = 0;
assign rom[2][11] = 0;
assign rom[2][12] = 0;
assign rom[2][13] = 0;
assign rom[2][14] = 0;
assign rom[2][15] = 0;
assign rom[2][16] = 0;
assign rom[2][17] = 0;
assign rom[2][18] = 0;
assign rom[2][19] = 0;
assign rom[2][20] = 0;
assign rom[2][21] = 0;
assign rom[2][22] = 0;
assign rom[2][23] = 0;
assign rom[2][24] = 0;
assign rom[2][25] = 0;
assign rom[2][26] = 0;
assign rom[2][27] = 0;
assign rom[3][0] = 0;
assign rom[3][1] = 0;
assign rom[3][2] = 0;
assign rom[3][3] = 0;
assign rom[3][4] = 0;
assign rom[3][5] = 0;
assign rom[3][6] = 0;
assign rom[3][7] = 0;
assign rom[3][8] = 0;
assign rom[3][9] = 0;
assign rom[3][10] = 116;
assign rom[3][11] = 125;
assign rom[3][12] = 171;
assign rom[3][13] = 255;
assign rom[3][14] = 255;
assign rom[3][15] = 150;
assign rom[3][16] = 93;
assign rom[3][17] = 0;
assign rom[3][18] = 0;
assign rom[3][19] = 0;
assign rom[3][20] = 0;
assign rom[3][21] = 0;
assign rom[3][22] = 0;
assign rom[3][23] = 0;
assign rom[3][24] = 0;
assign rom[3][25] = 0;
assign rom[3][26] = 0;
assign rom[3][27] = 0;
assign rom[4][0] = 0;
assign rom[4][1] = 0;
assign rom[4][2] = 0;
assign rom[4][3] = 0;
assign rom[4][4] = 0;
assign rom[4][5] = 0;
assign rom[4][6] = 0;
assign rom[4][7] = 0;
assign rom[4][8] = 0;
assign rom[4][9] = 169;
assign rom[4][10] = 253;
assign rom[4][11] = 253;
assign rom[4][12] = 253;
assign rom[4][13] = 253;
assign rom[4][14] = 253;
assign rom[4][15] = 253;
assign rom[4][16] = 218;
assign rom[4][17] = 30;
assign rom[4][18] = 0;
assign rom[4][19] = 0;
assign rom[4][20] = 0;
assign rom[4][21] = 0;
assign rom[4][22] = 0;
assign rom[4][23] = 0;
assign rom[4][24] = 0;
assign rom[4][25] = 0;
assign rom[4][26] = 0;
assign rom[4][27] = 0;
assign rom[5][0] = 0;
assign rom[5][1] = 0;
assign rom[5][2] = 0;
assign rom[5][3] = 0;
assign rom[5][4] = 0;
assign rom[5][5] = 0;
assign rom[5][6] = 0;
assign rom[5][7] = 0;
assign rom[5][8] = 169;
assign rom[5][9] = 253;
assign rom[5][10] = 253;
assign rom[5][11] = 253;
assign rom[5][12] = 213;
assign rom[5][13] = 142;
assign rom[5][14] = 176;
assign rom[5][15] = 253;
assign rom[5][16] = 253;
assign rom[5][17] = 122;
assign rom[5][18] = 0;
assign rom[5][19] = 0;
assign rom[5][20] = 0;
assign rom[5][21] = 0;
assign rom[5][22] = 0;
assign rom[5][23] = 0;
assign rom[5][24] = 0;
assign rom[5][25] = 0;
assign rom[5][26] = 0;
assign rom[5][27] = 0;
assign rom[6][0] = 0;
assign rom[6][1] = 0;
assign rom[6][2] = 0;
assign rom[6][3] = 0;
assign rom[6][4] = 0;
assign rom[6][5] = 0;
assign rom[6][6] = 0;
assign rom[6][7] = 52;
assign rom[6][8] = 250;
assign rom[6][9] = 253;
assign rom[6][10] = 210;
assign rom[6][11] = 32;
assign rom[6][12] = 12;
assign rom[6][13] = 0;
assign rom[6][14] = 6;
assign rom[6][15] = 206;
assign rom[6][16] = 253;
assign rom[6][17] = 140;
assign rom[6][18] = 0;
assign rom[6][19] = 0;
assign rom[6][20] = 0;
assign rom[6][21] = 0;
assign rom[6][22] = 0;
assign rom[6][23] = 0;
assign rom[6][24] = 0;
assign rom[6][25] = 0;
assign rom[6][26] = 0;
assign rom[6][27] = 0;
assign rom[7][0] = 0;
assign rom[7][1] = 0;
assign rom[7][2] = 0;
assign rom[7][3] = 0;
assign rom[7][4] = 0;
assign rom[7][5] = 0;
assign rom[7][6] = 0;
assign rom[7][7] = 77;
assign rom[7][8] = 251;
assign rom[7][9] = 210;
assign rom[7][10] = 25;
assign rom[7][11] = 0;
assign rom[7][12] = 0;
assign rom[7][13] = 0;
assign rom[7][14] = 122;
assign rom[7][15] = 248;
assign rom[7][16] = 253;
assign rom[7][17] = 65;
assign rom[7][18] = 0;
assign rom[7][19] = 0;
assign rom[7][20] = 0;
assign rom[7][21] = 0;
assign rom[7][22] = 0;
assign rom[7][23] = 0;
assign rom[7][24] = 0;
assign rom[7][25] = 0;
assign rom[7][26] = 0;
assign rom[7][27] = 0;
assign rom[8][0] = 0;
assign rom[8][1] = 0;
assign rom[8][2] = 0;
assign rom[8][3] = 0;
assign rom[8][4] = 0;
assign rom[8][5] = 0;
assign rom[8][6] = 0;
assign rom[8][7] = 0;
assign rom[8][8] = 31;
assign rom[8][9] = 18;
assign rom[8][10] = 0;
assign rom[8][11] = 0;
assign rom[8][12] = 0;
assign rom[8][13] = 0;
assign rom[8][14] = 209;
assign rom[8][15] = 253;
assign rom[8][16] = 253;
assign rom[8][17] = 65;
assign rom[8][18] = 0;
assign rom[8][19] = 0;
assign rom[8][20] = 0;
assign rom[8][21] = 0;
assign rom[8][22] = 0;
assign rom[8][23] = 0;
assign rom[8][24] = 0;
assign rom[8][25] = 0;
assign rom[8][26] = 0;
assign rom[8][27] = 0;
assign rom[9][0] = 0;
assign rom[9][1] = 0;
assign rom[9][2] = 0;
assign rom[9][3] = 0;
assign rom[9][4] = 0;
assign rom[9][5] = 0;
assign rom[9][6] = 0;
assign rom[9][7] = 0;
assign rom[9][8] = 0;
assign rom[9][9] = 0;
assign rom[9][10] = 0;
assign rom[9][11] = 0;
assign rom[9][12] = 0;
assign rom[9][13] = 117;
assign rom[9][14] = 247;
assign rom[9][15] = 253;
assign rom[9][16] = 198;
assign rom[9][17] = 10;
assign rom[9][18] = 0;
assign rom[9][19] = 0;
assign rom[9][20] = 0;
assign rom[9][21] = 0;
assign rom[9][22] = 0;
assign rom[9][23] = 0;
assign rom[9][24] = 0;
assign rom[9][25] = 0;
assign rom[9][26] = 0;
assign rom[9][27] = 0;
assign rom[10][0] = 0;
assign rom[10][1] = 0;
assign rom[10][2] = 0;
assign rom[10][3] = 0;
assign rom[10][4] = 0;
assign rom[10][5] = 0;
assign rom[10][6] = 0;
assign rom[10][7] = 0;
assign rom[10][8] = 0;
assign rom[10][9] = 0;
assign rom[10][10] = 0;
assign rom[10][11] = 0;
assign rom[10][12] = 76;
assign rom[10][13] = 247;
assign rom[10][14] = 253;
assign rom[10][15] = 231;
assign rom[10][16] = 63;
assign rom[10][17] = 0;
assign rom[10][18] = 0;
assign rom[10][19] = 0;
assign rom[10][20] = 0;
assign rom[10][21] = 0;
assign rom[10][22] = 0;
assign rom[10][23] = 0;
assign rom[10][24] = 0;
assign rom[10][25] = 0;
assign rom[10][26] = 0;
assign rom[10][27] = 0;
assign rom[11][0] = 0;
assign rom[11][1] = 0;
assign rom[11][2] = 0;
assign rom[11][3] = 0;
assign rom[11][4] = 0;
assign rom[11][5] = 0;
assign rom[11][6] = 0;
assign rom[11][7] = 0;
assign rom[11][8] = 0;
assign rom[11][9] = 0;
assign rom[11][10] = 0;
assign rom[11][11] = 0;
assign rom[11][12] = 128;
assign rom[11][13] = 253;
assign rom[11][14] = 253;
assign rom[11][15] = 144;
assign rom[11][16] = 0;
assign rom[11][17] = 0;
assign rom[11][18] = 0;
assign rom[11][19] = 0;
assign rom[11][20] = 0;
assign rom[11][21] = 0;
assign rom[11][22] = 0;
assign rom[11][23] = 0;
assign rom[11][24] = 0;
assign rom[11][25] = 0;
assign rom[11][26] = 0;
assign rom[11][27] = 0;
assign rom[12][0] = 0;
assign rom[12][1] = 0;
assign rom[12][2] = 0;
assign rom[12][3] = 0;
assign rom[12][4] = 0;
assign rom[12][5] = 0;
assign rom[12][6] = 0;
assign rom[12][7] = 0;
assign rom[12][8] = 0;
assign rom[12][9] = 0;
assign rom[12][10] = 0;
assign rom[12][11] = 176;
assign rom[12][12] = 246;
assign rom[12][13] = 253;
assign rom[12][14] = 159;
assign rom[12][15] = 12;
assign rom[12][16] = 0;
assign rom[12][17] = 0;
assign rom[12][18] = 0;
assign rom[12][19] = 0;
assign rom[12][20] = 0;
assign rom[12][21] = 0;
assign rom[12][22] = 0;
assign rom[12][23] = 0;
assign rom[12][24] = 0;
assign rom[12][25] = 0;
assign rom[12][26] = 0;
assign rom[12][27] = 0;
assign rom[13][0] = 0;
assign rom[13][1] = 0;
assign rom[13][2] = 0;
assign rom[13][3] = 0;
assign rom[13][4] = 0;
assign rom[13][5] = 0;
assign rom[13][6] = 0;
assign rom[13][7] = 0;
assign rom[13][8] = 0;
assign rom[13][9] = 0;
assign rom[13][10] = 25;
assign rom[13][11] = 234;
assign rom[13][12] = 253;
assign rom[13][13] = 233;
assign rom[13][14] = 35;
assign rom[13][15] = 0;
assign rom[13][16] = 0;
assign rom[13][17] = 0;
assign rom[13][18] = 0;
assign rom[13][19] = 0;
assign rom[13][20] = 0;
assign rom[13][21] = 0;
assign rom[13][22] = 0;
assign rom[13][23] = 0;
assign rom[13][24] = 0;
assign rom[13][25] = 0;
assign rom[13][26] = 0;
assign rom[13][27] = 0;
assign rom[14][0] = 0;
assign rom[14][1] = 0;
assign rom[14][2] = 0;
assign rom[14][3] = 0;
assign rom[14][4] = 0;
assign rom[14][5] = 0;
assign rom[14][6] = 0;
assign rom[14][7] = 0;
assign rom[14][8] = 0;
assign rom[14][9] = 0;
assign rom[14][10] = 198;
assign rom[14][11] = 253;
assign rom[14][12] = 253;
assign rom[14][13] = 141;
assign rom[14][14] = 0;
assign rom[14][15] = 0;
assign rom[14][16] = 0;
assign rom[14][17] = 0;
assign rom[14][18] = 0;
assign rom[14][19] = 0;
assign rom[14][20] = 0;
assign rom[14][21] = 0;
assign rom[14][22] = 0;
assign rom[14][23] = 0;
assign rom[14][24] = 0;
assign rom[14][25] = 0;
assign rom[14][26] = 0;
assign rom[14][27] = 0;
assign rom[15][0] = 0;
assign rom[15][1] = 0;
assign rom[15][2] = 0;
assign rom[15][3] = 0;
assign rom[15][4] = 0;
assign rom[15][5] = 0;
assign rom[15][6] = 0;
assign rom[15][7] = 0;
assign rom[15][8] = 0;
assign rom[15][9] = 78;
assign rom[15][10] = 248;
assign rom[15][11] = 253;
assign rom[15][12] = 189;
assign rom[15][13] = 12;
assign rom[15][14] = 0;
assign rom[15][15] = 0;
assign rom[15][16] = 0;
assign rom[15][17] = 0;
assign rom[15][18] = 0;
assign rom[15][19] = 0;
assign rom[15][20] = 0;
assign rom[15][21] = 0;
assign rom[15][22] = 0;
assign rom[15][23] = 0;
assign rom[15][24] = 0;
assign rom[15][25] = 0;
assign rom[15][26] = 0;
assign rom[15][27] = 0;
assign rom[16][0] = 0;
assign rom[16][1] = 0;
assign rom[16][2] = 0;
assign rom[16][3] = 0;
assign rom[16][4] = 0;
assign rom[16][5] = 0;
assign rom[16][6] = 0;
assign rom[16][7] = 0;
assign rom[16][8] = 19;
assign rom[16][9] = 200;
assign rom[16][10] = 253;
assign rom[16][11] = 253;
assign rom[16][12] = 141;
assign rom[16][13] = 0;
assign rom[16][14] = 0;
assign rom[16][15] = 0;
assign rom[16][16] = 0;
assign rom[16][17] = 0;
assign rom[16][18] = 0;
assign rom[16][19] = 0;
assign rom[16][20] = 0;
assign rom[16][21] = 0;
assign rom[16][22] = 0;
assign rom[16][23] = 0;
assign rom[16][24] = 0;
assign rom[16][25] = 0;
assign rom[16][26] = 0;
assign rom[16][27] = 0;
assign rom[17][0] = 0;
assign rom[17][1] = 0;
assign rom[17][2] = 0;
assign rom[17][3] = 0;
assign rom[17][4] = 0;
assign rom[17][5] = 0;
assign rom[17][6] = 0;
assign rom[17][7] = 0;
assign rom[17][8] = 134;
assign rom[17][9] = 253;
assign rom[17][10] = 253;
assign rom[17][11] = 173;
assign rom[17][12] = 12;
assign rom[17][13] = 0;
assign rom[17][14] = 0;
assign rom[17][15] = 0;
assign rom[17][16] = 0;
assign rom[17][17] = 0;
assign rom[17][18] = 0;
assign rom[17][19] = 0;
assign rom[17][20] = 0;
assign rom[17][21] = 0;
assign rom[17][22] = 0;
assign rom[17][23] = 0;
assign rom[17][24] = 0;
assign rom[17][25] = 0;
assign rom[17][26] = 0;
assign rom[17][27] = 0;
assign rom[18][0] = 0;
assign rom[18][1] = 0;
assign rom[18][2] = 0;
assign rom[18][3] = 0;
assign rom[18][4] = 0;
assign rom[18][5] = 0;
assign rom[18][6] = 0;
assign rom[18][7] = 0;
assign rom[18][8] = 248;
assign rom[18][9] = 253;
assign rom[18][10] = 253;
assign rom[18][11] = 25;
assign rom[18][12] = 0;
assign rom[18][13] = 0;
assign rom[18][14] = 0;
assign rom[18][15] = 0;
assign rom[18][16] = 0;
assign rom[18][17] = 0;
assign rom[18][18] = 0;
assign rom[18][19] = 0;
assign rom[18][20] = 0;
assign rom[18][21] = 0;
assign rom[18][22] = 0;
assign rom[18][23] = 0;
assign rom[18][24] = 0;
assign rom[18][25] = 0;
assign rom[18][26] = 0;
assign rom[18][27] = 0;
assign rom[19][0] = 0;
assign rom[19][1] = 0;
assign rom[19][2] = 0;
assign rom[19][3] = 0;
assign rom[19][4] = 0;
assign rom[19][5] = 0;
assign rom[19][6] = 0;
assign rom[19][7] = 0;
assign rom[19][8] = 248;
assign rom[19][9] = 253;
assign rom[19][10] = 253;
assign rom[19][11] = 43;
assign rom[19][12] = 20;
assign rom[19][13] = 20;
assign rom[19][14] = 20;
assign rom[19][15] = 20;
assign rom[19][16] = 5;
assign rom[19][17] = 0;
assign rom[19][18] = 5;
assign rom[19][19] = 20;
assign rom[19][20] = 20;
assign rom[19][21] = 37;
assign rom[19][22] = 150;
assign rom[19][23] = 150;
assign rom[19][24] = 150;
assign rom[19][25] = 147;
assign rom[19][26] = 10;
assign rom[19][27] = 0;
assign rom[20][0] = 0;
assign rom[20][1] = 0;
assign rom[20][2] = 0;
assign rom[20][3] = 0;
assign rom[20][4] = 0;
assign rom[20][5] = 0;
assign rom[20][6] = 0;
assign rom[20][7] = 0;
assign rom[20][8] = 248;
assign rom[20][9] = 253;
assign rom[20][10] = 253;
assign rom[20][11] = 253;
assign rom[20][12] = 253;
assign rom[20][13] = 253;
assign rom[20][14] = 253;
assign rom[20][15] = 253;
assign rom[20][16] = 168;
assign rom[20][17] = 143;
assign rom[20][18] = 166;
assign rom[20][19] = 253;
assign rom[20][20] = 253;
assign rom[20][21] = 253;
assign rom[20][22] = 253;
assign rom[20][23] = 253;
assign rom[20][24] = 253;
assign rom[20][25] = 253;
assign rom[20][26] = 123;
assign rom[20][27] = 0;
assign rom[21][0] = 0;
assign rom[21][1] = 0;
assign rom[21][2] = 0;
assign rom[21][3] = 0;
assign rom[21][4] = 0;
assign rom[21][5] = 0;
assign rom[21][6] = 0;
assign rom[21][7] = 0;
assign rom[21][8] = 174;
assign rom[21][9] = 253;
assign rom[21][10] = 253;
assign rom[21][11] = 253;
assign rom[21][12] = 253;
assign rom[21][13] = 253;
assign rom[21][14] = 253;
assign rom[21][15] = 253;
assign rom[21][16] = 253;
assign rom[21][17] = 253;
assign rom[21][18] = 253;
assign rom[21][19] = 253;
assign rom[21][20] = 249;
assign rom[21][21] = 247;
assign rom[21][22] = 247;
assign rom[21][23] = 169;
assign rom[21][24] = 117;
assign rom[21][25] = 117;
assign rom[21][26] = 57;
assign rom[21][27] = 0;
assign rom[22][0] = 0;
assign rom[22][1] = 0;
assign rom[22][2] = 0;
assign rom[22][3] = 0;
assign rom[22][4] = 0;
assign rom[22][5] = 0;
assign rom[22][6] = 0;
assign rom[22][7] = 0;
assign rom[22][8] = 0;
assign rom[22][9] = 118;
assign rom[22][10] = 123;
assign rom[22][11] = 123;
assign rom[22][12] = 123;
assign rom[22][13] = 166;
assign rom[22][14] = 253;
assign rom[22][15] = 253;
assign rom[22][16] = 253;
assign rom[22][17] = 155;
assign rom[22][18] = 123;
assign rom[22][19] = 123;
assign rom[22][20] = 41;
assign rom[22][21] = 0;
assign rom[22][22] = 0;
assign rom[22][23] = 0;
assign rom[22][24] = 0;
assign rom[22][25] = 0;
assign rom[22][26] = 0;
assign rom[22][27] = 0;
assign rom[23][0] = 0;
assign rom[23][1] = 0;
assign rom[23][2] = 0;
assign rom[23][3] = 0;
assign rom[23][4] = 0;
assign rom[23][5] = 0;
assign rom[23][6] = 0;
assign rom[23][7] = 0;
assign rom[23][8] = 0;
assign rom[23][9] = 0;
assign rom[23][10] = 0;
assign rom[23][11] = 0;
assign rom[23][12] = 0;
assign rom[23][13] = 0;
assign rom[23][14] = 0;
assign rom[23][15] = 0;
assign rom[23][16] = 0;
assign rom[23][17] = 0;
assign rom[23][18] = 0;
assign rom[23][19] = 0;
assign rom[23][20] = 0;
assign rom[23][21] = 0;
assign rom[23][22] = 0;
assign rom[23][23] = 0;
assign rom[23][24] = 0;
assign rom[23][25] = 0;
assign rom[23][26] = 0;
assign rom[23][27] = 0;
assign rom[24][0] = 0;
assign rom[24][1] = 0;
assign rom[24][2] = 0;
assign rom[24][3] = 0;
assign rom[24][4] = 0;
assign rom[24][5] = 0;
assign rom[24][6] = 0;
assign rom[24][7] = 0;
assign rom[24][8] = 0;
assign rom[24][9] = 0;
assign rom[24][10] = 0;
assign rom[24][11] = 0;
assign rom[24][12] = 0;
assign rom[24][13] = 0;
assign rom[24][14] = 0;
assign rom[24][15] = 0;
assign rom[24][16] = 0;
assign rom[24][17] = 0;
assign rom[24][18] = 0;
assign rom[24][19] = 0;
assign rom[24][20] = 0;
assign rom[24][21] = 0;
assign rom[24][22] = 0;
assign rom[24][23] = 0;
assign rom[24][24] = 0;
assign rom[24][25] = 0;
assign rom[24][26] = 0;
assign rom[24][27] = 0;
assign rom[25][0] = 0;
assign rom[25][1] = 0;
assign rom[25][2] = 0;
assign rom[25][3] = 0;
assign rom[25][4] = 0;
assign rom[25][5] = 0;
assign rom[25][6] = 0;
assign rom[25][7] = 0;
assign rom[25][8] = 0;
assign rom[25][9] = 0;
assign rom[25][10] = 0;
assign rom[25][11] = 0;
assign rom[25][12] = 0;
assign rom[25][13] = 0;
assign rom[25][14] = 0;
assign rom[25][15] = 0;
assign rom[25][16] = 0;
assign rom[25][17] = 0;
assign rom[25][18] = 0;
assign rom[25][19] = 0;
assign rom[25][20] = 0;
assign rom[25][21] = 0;
assign rom[25][22] = 0;
assign rom[25][23] = 0;
assign rom[25][24] = 0;
assign rom[25][25] = 0;
assign rom[25][26] = 0;
assign rom[25][27] = 0;
assign rom[26][0] = 0;
assign rom[26][1] = 0;
assign rom[26][2] = 0;
assign rom[26][3] = 0;
assign rom[26][4] = 0;
assign rom[26][5] = 0;
assign rom[26][6] = 0;
assign rom[26][7] = 0;
assign rom[26][8] = 0;
assign rom[26][9] = 0;
assign rom[26][10] = 0;
assign rom[26][11] = 0;
assign rom[26][12] = 0;
assign rom[26][13] = 0;
assign rom[26][14] = 0;
assign rom[26][15] = 0;
assign rom[26][16] = 0;
assign rom[26][17] = 0;
assign rom[26][18] = 0;
assign rom[26][19] = 0;
assign rom[26][20] = 0;
assign rom[26][21] = 0;
assign rom[26][22] = 0;
assign rom[26][23] = 0;
assign rom[26][24] = 0;
assign rom[26][25] = 0;
assign rom[26][26] = 0;
assign rom[26][27] = 0;
assign rom[27][0] = 0;
assign rom[27][1] = 0;
assign rom[27][2] = 0;
assign rom[27][3] = 0;
assign rom[27][4] = 0;
assign rom[27][5] = 0;
assign rom[27][6] = 0;
assign rom[27][7] = 0;
assign rom[27][8] = 0;
assign rom[27][9] = 0;
assign rom[27][10] = 0;
assign rom[27][11] = 0;
assign rom[27][12] = 0;
assign rom[27][13] = 0;
assign rom[27][14] = 0;
assign rom[27][15] = 0;
assign rom[27][16] = 0;
assign rom[27][17] = 0;
assign rom[27][18] = 0;
assign rom[27][19] = 0;
assign rom[27][20] = 0;
assign rom[27][21] = 0;
assign rom[27][22] = 0;
assign rom[27][23] = 0;
assign rom[27][24] = 0;
assign rom[27][25] = 0;
assign rom[27][26] = 0;
assign rom[27][27] = 0;


endmodule