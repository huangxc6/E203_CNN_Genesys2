/******************************************************************************
*
*  Authors:   Chengyi Zhang
*     Date:   2023/4/20
*   Method:   
*  Version:   
*  Content:  
* 
******************************************************************************/

module conv_weight_buffer (
    output             [   7: 0]        o_weight [ 8:0]             ,
    output             [   7: 0]        o_bias 
);

logic   [   7: 0]   rom    [   8: 0];

assign o_weight = rom;
assign o_bias   = 19;

// # conv_0_filter_0
// 20 60 18 56 88 105 40 74 101

assign rom[0] = 20  ;
assign rom[1] = 60  ;
assign rom[2] = 18  ;
assign rom[3] = 56  ;
assign rom[4] = 88  ;
assign rom[5] = 105 ;
assign rom[6] = 40  ;
assign rom[7] = 74  ;
assign rom[8] = 101 ;

endmodule

module fc_weight_buffer (
    input              [   4: 0]        i_addr                     ,
    output             [   7: 0]        o_weight      [25:0][9:0]  ,
    output             [   7: 0]        o_bias              [9:0]              
);

logic   [   7: 0]   rom    [   675: 0][   9: 0];

generate
    for (genvar i = 0; i < 26; i++) begin
        for (genvar j = 0; j < 10; j++) begin
            assign o_weight[i][j] = rom[26*i_addr+i][j];
        end
    end
endgenerate

// -4 15 -3 -8 5 10 -2 9 -18 -3

assign o_bias[0] = -4 ;
assign o_bias[1] = 15 ;
assign o_bias[2] = -3 ;
assign o_bias[3] = -8 ;
assign o_bias[4] = 5  ;
assign o_bias[5] = 10 ;
assign o_bias[6] = -2 ;
assign o_bias[7] = 9  ;
assign o_bias[8] = -18;
assign o_bias[9] = -3 ;

assign rom[0][0] = -7;
assign rom[0][1] = 29;
assign rom[0][2] = -5;
assign rom[0][3] = -10;
assign rom[0][4] = 6;
assign rom[0][5] = 10;
assign rom[0][6] = 5;
assign rom[0][7] = 16;
assign rom[0][8] = -29;
assign rom[0][9] = 4;
assign rom[1][0] = 1;
assign rom[1][1] = 27;
assign rom[1][2] = -6;
assign rom[1][3] = -16;
assign rom[1][4] = 10;
assign rom[1][5] = 23;
assign rom[1][6] = 1;
assign rom[1][7] = 8;
assign rom[1][8] = -20;
assign rom[1][9] = -8;
assign rom[2][0] = 1;
assign rom[2][1] = 16;
assign rom[2][2] = -9;
assign rom[2][3] = -12;
assign rom[2][4] = 9;
assign rom[2][5] = 7;
assign rom[2][6] = -8;
assign rom[2][7] = 10;
assign rom[2][8] = -26;
assign rom[2][9] = 2;
assign rom[3][0] = -15;
assign rom[3][1] = 26;
assign rom[3][2] = -9;
assign rom[3][3] = -15;
assign rom[3][4] = 1;
assign rom[3][5] = 9;
assign rom[3][6] = -1;
assign rom[3][7] = 8;
assign rom[3][8] = -15;
assign rom[3][9] = 1;
assign rom[4][0] = -14;
assign rom[4][1] = 30;
assign rom[4][2] = -4;
assign rom[4][3] = -11;
assign rom[4][4] = 13;
assign rom[4][5] = 18;
assign rom[4][6] = 3;
assign rom[4][7] = 13;
assign rom[4][8] = -18;
assign rom[4][9] = 0;
assign rom[5][0] = -2;
assign rom[5][1] = 23;
assign rom[5][2] = -5;
assign rom[5][3] = -20;
assign rom[5][4] = 3;
assign rom[5][5] = 8;
assign rom[5][6] = 8;
assign rom[5][7] = 13;
assign rom[5][8] = -21;
assign rom[5][9] = -14;
assign rom[6][0] = -14;
assign rom[6][1] = 19;
assign rom[6][2] = 1;
assign rom[6][3] = -11;
assign rom[6][4] = -3;
assign rom[6][5] = 22;
assign rom[6][6] = 10;
assign rom[6][7] = 2;
assign rom[6][8] = -27;
assign rom[6][9] = 0;
assign rom[7][0] = -11;
assign rom[7][1] = 14;
assign rom[7][2] = -6;
assign rom[7][3] = -16;
assign rom[7][4] = -3;
assign rom[7][5] = 6;
assign rom[7][6] = 19;
assign rom[7][7] = 4;
assign rom[7][8] = -25;
assign rom[7][9] = -11;
assign rom[8][0] = -17;
assign rom[8][1] = 17;
assign rom[8][2] = -4;
assign rom[8][3] = -20;
assign rom[8][4] = -4;
assign rom[8][5] = 11;
assign rom[8][6] = 12;
assign rom[8][7] = 14;
assign rom[8][8] = -22;
assign rom[8][9] = -11;
assign rom[9][0] = -19;
assign rom[9][1] = 25;
assign rom[9][2] = -14;
assign rom[9][3] = -13;
assign rom[9][4] = -19;
assign rom[9][5] = 1;
assign rom[9][6] = 25;
assign rom[9][7] = 11;
assign rom[9][8] = -20;
assign rom[9][9] = -8;
assign rom[10][0] = -11;
assign rom[10][1] = 14;
assign rom[10][2] = -13;
assign rom[10][3] = -23;
assign rom[10][4] = -19;
assign rom[10][5] = 0;
assign rom[10][6] = 14;
assign rom[10][7] = 14;
assign rom[10][8] = -22;
assign rom[10][9] = -16;
assign rom[11][0] = -12;
assign rom[11][1] = 20;
assign rom[11][2] = 2;
assign rom[11][3] = -19;
assign rom[11][4] = -16;
assign rom[11][5] = -2;
assign rom[11][6] = 16;
assign rom[11][7] = 3;
assign rom[11][8] = -23;
assign rom[11][9] = -5;
assign rom[12][0] = -12;
assign rom[12][1] = 10;
assign rom[12][2] = -9;
assign rom[12][3] = -21;
assign rom[12][4] = -26;
assign rom[12][5] = 10;
assign rom[12][6] = 16;
assign rom[12][7] = -3;
assign rom[12][8] = -27;
assign rom[12][9] = -6;
assign rom[13][0] = -18;
assign rom[13][1] = 24;
assign rom[13][2] = -7;
assign rom[13][3] = -24;
assign rom[13][4] = -19;
assign rom[13][5] = -3;
assign rom[13][6] = 16;
assign rom[13][7] = 2;
assign rom[13][8] = -27;
assign rom[13][9] = -14;
assign rom[14][0] = -14;
assign rom[14][1] = 13;
assign rom[14][2] = -8;
assign rom[14][3] = -12;
assign rom[14][4] = -10;
assign rom[14][5] = 7;
assign rom[14][6] = 7;
assign rom[14][7] = 3;
assign rom[14][8] = -30;
assign rom[14][9] = -13;
assign rom[15][0] = -13;
assign rom[15][1] = 7;
assign rom[15][2] = -3;
assign rom[15][3] = -25;
assign rom[15][4] = -11;
assign rom[15][5] = 5;
assign rom[15][6] = 6;
assign rom[15][7] = 8;
assign rom[15][8] = -32;
assign rom[15][9] = -2;
assign rom[16][0] = -7;
assign rom[16][1] = 10;
assign rom[16][2] = -3;
assign rom[16][3] = -13;
assign rom[16][4] = -11;
assign rom[16][5] = -2;
assign rom[16][6] = 17;
assign rom[16][7] = -1;
assign rom[16][8] = -33;
assign rom[16][9] = -10;
assign rom[17][0] = -12;
assign rom[17][1] = 0;
assign rom[17][2] = -8;
assign rom[17][3] = -29;
assign rom[17][4] = -3;
assign rom[17][5] = 12;
assign rom[17][6] = 24;
assign rom[17][7] = 10;
assign rom[17][8] = -34;
assign rom[17][9] = -8;
assign rom[18][0] = -14;
assign rom[18][1] = 12;
assign rom[18][2] = -17;
assign rom[18][3] = -14;
assign rom[18][4] = -1;
assign rom[18][5] = 6;
assign rom[18][6] = 15;
assign rom[18][7] = 12;
assign rom[18][8] = -21;
assign rom[18][9] = -3;
assign rom[19][0] = -17;
assign rom[19][1] = 18;
assign rom[19][2] = -19;
assign rom[19][3] = -24;
assign rom[19][4] = 8;
assign rom[19][5] = 9;
assign rom[19][6] = 19;
assign rom[19][7] = 16;
assign rom[19][8] = -23;
assign rom[19][9] = -14;
assign rom[20][0] = -11;
assign rom[20][1] = 21;
assign rom[20][2] = -2;
assign rom[20][3] = -10;
assign rom[20][4] = -7;
assign rom[20][5] = 10;
assign rom[20][6] = 4;
assign rom[20][7] = 15;
assign rom[20][8] = -32;
assign rom[20][9] = -8;
assign rom[21][0] = -11;
assign rom[21][1] = 19;
assign rom[21][2] = -11;
assign rom[21][3] = -19;
assign rom[21][4] = 5;
assign rom[21][5] = 12;
assign rom[21][6] = 0;
assign rom[21][7] = 6;
assign rom[21][8] = -19;
assign rom[21][9] = -4;
assign rom[22][0] = -3;
assign rom[22][1] = 19;
assign rom[22][2] = -12;
assign rom[22][3] = -16;
assign rom[22][4] = 15;
assign rom[22][5] = 6;
assign rom[22][6] = 10;
assign rom[22][7] = 7;
assign rom[22][8] = -25;
assign rom[22][9] = -7;
assign rom[23][0] = -6;
assign rom[23][1] = 16;
assign rom[23][2] = -7;
assign rom[23][3] = -21;
assign rom[23][4] = -1;
assign rom[23][5] = 20;
assign rom[23][6] = 0;
assign rom[23][7] = 10;
assign rom[23][8] = -15;
assign rom[23][9] = 3;
assign rom[24][0] = -3;
assign rom[24][1] = 16;
assign rom[24][2] = -6;
assign rom[24][3] = -16;
assign rom[24][4] = 6;
assign rom[24][5] = 23;
assign rom[24][6] = 3;
assign rom[24][7] = 6;
assign rom[24][8] = -29;
assign rom[24][9] = -11;
assign rom[25][0] = -1;
assign rom[25][1] = 20;
assign rom[25][2] = -8;
assign rom[25][3] = -4;
assign rom[25][4] = 2;
assign rom[25][5] = 19;
assign rom[25][6] = 3;
assign rom[25][7] = 19;
assign rom[25][8] = -15;
assign rom[25][9] = 0;
assign rom[26][0] = -2;
assign rom[26][1] = 18;
assign rom[26][2] = -7;
assign rom[26][3] = -21;
assign rom[26][4] = 14;
assign rom[26][5] = 21;
assign rom[26][6] = 5;
assign rom[26][7] = 20;
assign rom[26][8] = -26;
assign rom[26][9] = -6;
assign rom[27][0] = -11;
assign rom[27][1] = 32;
assign rom[27][2] = -12;
assign rom[27][3] = -14;
assign rom[27][4] = 6;
assign rom[27][5] = 6;
assign rom[27][6] = 2;
assign rom[27][7] = 11;
assign rom[27][8] = -23;
assign rom[27][9] = -11;
assign rom[28][0] = -12;
assign rom[28][1] = 28;
assign rom[28][2] = -4;
assign rom[28][3] = -14;
assign rom[28][4] = 1;
assign rom[28][5] = 23;
assign rom[28][6] = -10;
assign rom[28][7] = 14;
assign rom[28][8] = -28;
assign rom[28][9] = -9;
assign rom[29][0] = -15;
assign rom[29][1] = 20;
assign rom[29][2] = -4;
assign rom[29][3] = -6;
assign rom[29][4] = 8;
assign rom[29][5] = 12;
assign rom[29][6] = 2;
assign rom[29][7] = 13;
assign rom[29][8] = -33;
assign rom[29][9] = -13;
assign rom[30][0] = 1;
assign rom[30][1] = 16;
assign rom[30][2] = -13;
assign rom[30][3] = -19;
assign rom[30][4] = 9;
assign rom[30][5] = 7;
assign rom[30][6] = 3;
assign rom[30][7] = 8;
assign rom[30][8] = -19;
assign rom[30][9] = -11;
assign rom[31][0] = -2;
assign rom[31][1] = 21;
assign rom[31][2] = -1;
assign rom[31][3] = -6;
assign rom[31][4] = 2;
assign rom[31][5] = 14;
assign rom[31][6] = 10;
assign rom[31][7] = 4;
assign rom[31][8] = -34;
assign rom[31][9] = 0;
assign rom[32][0] = -8;
assign rom[32][1] = 8;
assign rom[32][2] = -8;
assign rom[32][3] = -7;
assign rom[32][4] = -14;
assign rom[32][5] = 6;
assign rom[32][6] = 22;
assign rom[32][7] = 2;
assign rom[32][8] = -18;
assign rom[32][9] = -7;
assign rom[33][0] = -21;
assign rom[33][1] = -1;
assign rom[33][2] = 10;
assign rom[33][3] = -15;
assign rom[33][4] = -9;
assign rom[33][5] = 14;
assign rom[33][6] = 23;
assign rom[33][7] = 4;
assign rom[33][8] = -18;
assign rom[33][9] = -13;
assign rom[34][0] = -24;
assign rom[34][1] = -2;
assign rom[34][2] = 7;
assign rom[34][3] = -1;
assign rom[34][4] = -26;
assign rom[34][5] = 1;
assign rom[34][6] = 21;
assign rom[34][7] = 8;
assign rom[34][8] = -21;
assign rom[34][9] = -6;
assign rom[35][0] = -14;
assign rom[35][1] = -1;
assign rom[35][2] = 5;
assign rom[35][3] = 5;
assign rom[35][4] = -29;
assign rom[35][5] = -1;
assign rom[35][6] = 28;
assign rom[35][7] = 8;
assign rom[35][8] = -25;
assign rom[35][9] = -9;
assign rom[36][0] = -25;
assign rom[36][1] = -10;
assign rom[36][2] = 15;
assign rom[36][3] = -1;
assign rom[36][4] = -43;
assign rom[36][5] = -3;
assign rom[36][6] = 31;
assign rom[36][7] = -6;
assign rom[36][8] = -38;
assign rom[36][9] = -19;
assign rom[37][0] = -12;
assign rom[37][1] = -11;
assign rom[37][2] = 12;
assign rom[37][3] = 15;
assign rom[37][4] = -40;
assign rom[37][5] = -3;
assign rom[37][6] = 30;
assign rom[37][7] = 7;
assign rom[37][8] = -30;
assign rom[37][9] = -9;
assign rom[38][0] = -23;
assign rom[38][1] = -3;
assign rom[38][2] = 3;
assign rom[38][3] = 7;
assign rom[38][4] = -46;
assign rom[38][5] = -9;
assign rom[38][6] = 27;
assign rom[38][7] = 3;
assign rom[38][8] = -25;
assign rom[38][9] = -11;
assign rom[39][0] = -19;
assign rom[39][1] = -1;
assign rom[39][2] = -4;
assign rom[39][3] = 17;
assign rom[39][4] = -46;
assign rom[39][5] = -6;
assign rom[39][6] = 15;
assign rom[39][7] = 1;
assign rom[39][8] = -35;
assign rom[39][9] = -15;
assign rom[40][0] = -28;
assign rom[40][1] = 7;
assign rom[40][2] = -4;
assign rom[40][3] = 14;
assign rom[40][4] = -23;
assign rom[40][5] = -12;
assign rom[40][6] = 15;
assign rom[40][7] = 1;
assign rom[40][8] = -24;
assign rom[40][9] = -20;
assign rom[41][0] = -25;
assign rom[41][1] = -2;
assign rom[41][2] = -2;
assign rom[41][3] = 13;
assign rom[41][4] = -19;
assign rom[41][5] = 0;
assign rom[41][6] = 17;
assign rom[41][7] = 3;
assign rom[41][8] = -30;
assign rom[41][9] = -8;
assign rom[42][0] = -26;
assign rom[42][1] = -23;
assign rom[42][2] = -5;
assign rom[42][3] = 6;
assign rom[42][4] = -26;
assign rom[42][5] = -3;
assign rom[42][6] = 25;
assign rom[42][7] = 4;
assign rom[42][8] = -36;
assign rom[42][9] = -17;
assign rom[43][0] = -36;
assign rom[43][1] = -25;
assign rom[43][2] = -15;
assign rom[43][3] = -5;
assign rom[43][4] = -19;
assign rom[43][5] = -6;
assign rom[43][6] = 35;
assign rom[43][7] = -8;
assign rom[43][8] = -34;
assign rom[43][9] = -5;
assign rom[44][0] = -18;
assign rom[44][1] = -24;
assign rom[44][2] = -14;
assign rom[44][3] = 1;
assign rom[44][4] = -11;
assign rom[44][5] = -11;
assign rom[44][6] = 25;
assign rom[44][7] = 11;
assign rom[44][8] = -19;
assign rom[44][9] = -16;
assign rom[45][0] = -25;
assign rom[45][1] = -6;
assign rom[45][2] = -19;
assign rom[45][3] = -10;
assign rom[45][4] = -1;
assign rom[45][5] = 7;
assign rom[45][6] = 37;
assign rom[45][7] = 2;
assign rom[45][8] = -27;
assign rom[45][9] = -8;
assign rom[46][0] = -23;
assign rom[46][1] = -1;
assign rom[46][2] = -27;
assign rom[46][3] = -19;
assign rom[46][4] = -5;
assign rom[46][5] = 6;
assign rom[46][6] = 35;
assign rom[46][7] = 2;
assign rom[46][8] = -28;
assign rom[46][9] = -12;
assign rom[47][0] = -21;
assign rom[47][1] = 13;
assign rom[47][2] = -13;
assign rom[47][3] = -17;
assign rom[47][4] = -9;
assign rom[47][5] = -2;
assign rom[47][6] = 31;
assign rom[47][7] = 18;
assign rom[47][8] = -16;
assign rom[47][9] = 2;
assign rom[48][0] = -4;
assign rom[48][1] = 24;
assign rom[48][2] = -2;
assign rom[48][3] = -24;
assign rom[48][4] = 9;
assign rom[48][5] = 8;
assign rom[48][6] = 10;
assign rom[48][7] = 13;
assign rom[48][8] = -32;
assign rom[48][9] = -2;
assign rom[49][0] = -1;
assign rom[49][1] = 18;
assign rom[49][2] = -4;
assign rom[49][3] = -17;
assign rom[49][4] = 13;
assign rom[49][5] = 17;
assign rom[49][6] = 12;
assign rom[49][7] = 2;
assign rom[49][8] = -31;
assign rom[49][9] = -2;
assign rom[50][0] = -5;
assign rom[50][1] = 27;
assign rom[50][2] = -2;
assign rom[50][3] = -8;
assign rom[50][4] = 13;
assign rom[50][5] = 11;
assign rom[50][6] = -3;
assign rom[50][7] = 17;
assign rom[50][8] = -22;
assign rom[50][9] = 0;
assign rom[51][0] = -14;
assign rom[51][1] = 28;
assign rom[51][2] = -1;
assign rom[51][3] = -16;
assign rom[51][4] = 8;
assign rom[51][5] = 20;
assign rom[51][6] = 6;
assign rom[51][7] = 12;
assign rom[51][8] = -32;
assign rom[51][9] = 1;
assign rom[52][0] = -10;
assign rom[52][1] = 26;
assign rom[52][2] = -6;
assign rom[52][3] = -6;
assign rom[52][4] = 6;
assign rom[52][5] = 8;
assign rom[52][6] = -3;
assign rom[52][7] = 14;
assign rom[52][8] = -21;
assign rom[52][9] = 5;
assign rom[53][0] = -3;
assign rom[53][1] = 31;
assign rom[53][2] = -7;
assign rom[53][3] = -13;
assign rom[53][4] = 6;
assign rom[53][5] = 5;
assign rom[53][6] = -1;
assign rom[53][7] = 2;
assign rom[53][8] = -22;
assign rom[53][9] = -12;
assign rom[54][0] = -8;
assign rom[54][1] = 19;
assign rom[54][2] = 2;
assign rom[54][3] = -2;
assign rom[54][4] = -1;
assign rom[54][5] = 15;
assign rom[54][6] = -9;
assign rom[54][7] = 7;
assign rom[54][8] = -26;
assign rom[54][9] = -10;
assign rom[55][0] = -13;
assign rom[55][1] = 25;
assign rom[55][2] = -10;
assign rom[55][3] = 2;
assign rom[55][4] = 10;
assign rom[55][5] = 1;
assign rom[55][6] = 8;
assign rom[55][7] = 16;
assign rom[55][8] = -17;
assign rom[55][9] = -1;
assign rom[56][0] = -11;
assign rom[56][1] = 16;
assign rom[56][2] = -8;
assign rom[56][3] = 4;
assign rom[56][4] = -3;
assign rom[56][5] = 8;
assign rom[56][6] = -3;
assign rom[56][7] = 2;
assign rom[56][8] = -20;
assign rom[56][9] = -13;
assign rom[57][0] = -9;
assign rom[57][1] = 4;
assign rom[57][2] = -6;
assign rom[57][3] = 5;
assign rom[57][4] = -10;
assign rom[57][5] = 2;
assign rom[57][6] = 15;
assign rom[57][7] = -5;
assign rom[57][8] = -24;
assign rom[57][9] = -10;
assign rom[58][0] = -12;
assign rom[58][1] = -1;
assign rom[58][2] = 5;
assign rom[58][3] = 13;
assign rom[58][4] = -18;
assign rom[58][5] = -6;
assign rom[58][6] = 8;
assign rom[58][7] = -2;
assign rom[58][8] = -28;
assign rom[58][9] = -14;
assign rom[59][0] = -16;
assign rom[59][1] = -15;
assign rom[59][2] = 17;
assign rom[59][3] = 18;
assign rom[59][4] = -11;
assign rom[59][5] = -22;
assign rom[59][6] = 22;
assign rom[59][7] = -8;
assign rom[59][8] = -27;
assign rom[59][9] = -17;
assign rom[60][0] = -4;
assign rom[60][1] = -9;
assign rom[60][2] = 15;
assign rom[60][3] = 12;
assign rom[60][4] = -29;
assign rom[60][5] = -10;
assign rom[60][6] = 20;
assign rom[60][7] = -9;
assign rom[60][8] = -12;
assign rom[60][9] = -13;
assign rom[61][0] = -11;
assign rom[61][1] = -11;
assign rom[61][2] = 23;
assign rom[61][3] = 17;
assign rom[61][4] = -31;
assign rom[61][5] = -10;
assign rom[61][6] = 10;
assign rom[61][7] = -15;
assign rom[61][8] = -4;
assign rom[61][9] = -12;
assign rom[62][0] = -12;
assign rom[62][1] = 2;
assign rom[62][2] = 19;
assign rom[62][3] = 17;
assign rom[62][4] = -28;
assign rom[62][5] = -15;
assign rom[62][6] = 9;
assign rom[62][7] = -13;
assign rom[62][8] = -8;
assign rom[62][9] = -19;
assign rom[63][0] = -14;
assign rom[63][1] = -2;
assign rom[63][2] = 18;
assign rom[63][3] = 24;
assign rom[63][4] = -46;
assign rom[63][5] = -15;
assign rom[63][6] = 10;
assign rom[63][7] = -17;
assign rom[63][8] = -3;
assign rom[63][9] = -28;
assign rom[64][0] = -17;
assign rom[64][1] = -1;
assign rom[64][2] = 10;
assign rom[64][3] = 12;
assign rom[64][4] = -51;
assign rom[64][5] = -23;
assign rom[64][6] = 7;
assign rom[64][7] = -12;
assign rom[64][8] = 0;
assign rom[64][9] = -38;
assign rom[65][0] = -10;
assign rom[65][1] = 15;
assign rom[65][2] = 18;
assign rom[65][3] = 8;
assign rom[65][4] = -30;
assign rom[65][5] = -4;
assign rom[65][6] = 6;
assign rom[65][7] = -11;
assign rom[65][8] = 0;
assign rom[65][9] = -28;
assign rom[66][0] = -26;
assign rom[66][1] = 12;
assign rom[66][2] = 15;
assign rom[66][3] = 23;
assign rom[66][4] = -33;
assign rom[66][5] = 2;
assign rom[66][6] = 10;
assign rom[66][7] = -21;
assign rom[66][8] = -8;
assign rom[66][9] = -36;
assign rom[67][0] = -10;
assign rom[67][1] = -3;
assign rom[67][2] = 11;
assign rom[67][3] = 5;
assign rom[67][4] = -30;
assign rom[67][5] = 1;
assign rom[67][6] = 23;
assign rom[67][7] = -15;
assign rom[67][8] = -9;
assign rom[67][9] = -35;
assign rom[68][0] = -30;
assign rom[68][1] = -19;
assign rom[68][2] = -4;
assign rom[68][3] = 6;
assign rom[68][4] = -12;
assign rom[68][5] = -10;
assign rom[68][6] = 20;
assign rom[68][7] = -14;
assign rom[68][8] = -12;
assign rom[68][9] = -27;
assign rom[69][0] = -19;
assign rom[69][1] = -14;
assign rom[69][2] = -8;
assign rom[69][3] = 14;
assign rom[69][4] = -5;
assign rom[69][5] = -3;
assign rom[69][6] = 35;
assign rom[69][7] = -6;
assign rom[69][8] = -13;
assign rom[69][9] = -30;
assign rom[70][0] = -26;
assign rom[70][1] = -13;
assign rom[70][2] = -4;
assign rom[70][3] = -8;
assign rom[70][4] = -5;
assign rom[70][5] = 1;
assign rom[70][6] = 38;
assign rom[70][7] = -15;
assign rom[70][8] = -7;
assign rom[70][9] = -13;
assign rom[71][0] = -17;
assign rom[71][1] = -8;
assign rom[71][2] = -11;
assign rom[71][3] = -15;
assign rom[71][4] = 3;
assign rom[71][5] = -2;
assign rom[71][6] = 44;
assign rom[71][7] = -5;
assign rom[71][8] = -20;
assign rom[71][9] = -23;
assign rom[72][0] = -12;
assign rom[72][1] = 4;
assign rom[72][2] = -16;
assign rom[72][3] = -35;
assign rom[72][4] = 0;
assign rom[72][5] = -4;
assign rom[72][6] = 43;
assign rom[72][7] = 2;
assign rom[72][8] = -23;
assign rom[72][9] = -9;
assign rom[73][0] = -17;
assign rom[73][1] = 8;
assign rom[73][2] = -34;
assign rom[73][3] = -23;
assign rom[73][4] = 12;
assign rom[73][5] = 8;
assign rom[73][6] = 34;
assign rom[73][7] = 7;
assign rom[73][8] = -17;
assign rom[73][9] = -2;
assign rom[74][0] = -12;
assign rom[74][1] = 4;
assign rom[74][2] = -10;
assign rom[74][3] = -27;
assign rom[74][4] = 10;
assign rom[74][5] = 3;
assign rom[74][6] = 33;
assign rom[74][7] = 10;
assign rom[74][8] = -19;
assign rom[74][9] = -1;
assign rom[75][0] = -17;
assign rom[75][1] = 17;
assign rom[75][2] = -14;
assign rom[75][3] = -23;
assign rom[75][4] = 14;
assign rom[75][5] = 15;
assign rom[75][6] = 10;
assign rom[75][7] = 2;
assign rom[75][8] = -30;
assign rom[75][9] = 2;
assign rom[76][0] = -11;
assign rom[76][1] = 17;
assign rom[76][2] = 3;
assign rom[76][3] = -19;
assign rom[76][4] = 9;
assign rom[76][5] = 3;
assign rom[76][6] = -5;
assign rom[76][7] = 17;
assign rom[76][8] = -11;
assign rom[76][9] = -11;
assign rom[77][0] = -7;
assign rom[77][1] = 26;
assign rom[77][2] = -5;
assign rom[77][3] = -6;
assign rom[77][4] = 14;
assign rom[77][5] = 15;
assign rom[77][6] = -1;
assign rom[77][7] = 19;
assign rom[77][8] = -19;
assign rom[77][9] = 0;
assign rom[78][0] = -10;
assign rom[78][1] = 25;
assign rom[78][2] = 0;
assign rom[78][3] = -6;
assign rom[78][4] = 13;
assign rom[78][5] = 15;
assign rom[78][6] = 7;
assign rom[78][7] = 16;
assign rom[78][8] = -30;
assign rom[78][9] = 1;
assign rom[79][0] = -13;
assign rom[79][1] = 24;
assign rom[79][2] = -8;
assign rom[79][3] = -5;
assign rom[79][4] = 17;
assign rom[79][5] = 11;
assign rom[79][6] = -3;
assign rom[79][7] = 9;
assign rom[79][8] = -31;
assign rom[79][9] = 0;
assign rom[80][0] = -5;
assign rom[80][1] = 11;
assign rom[80][2] = -1;
assign rom[80][3] = -6;
assign rom[80][4] = 2;
assign rom[80][5] = 12;
assign rom[80][6] = -7;
assign rom[80][7] = 5;
assign rom[80][8] = -27;
assign rom[80][9] = -12;
assign rom[81][0] = -8;
assign rom[81][1] = 5;
assign rom[81][2] = -6;
assign rom[81][3] = 16;
assign rom[81][4] = 12;
assign rom[81][5] = -7;
assign rom[81][6] = -13;
assign rom[81][7] = 0;
assign rom[81][8] = -23;
assign rom[81][9] = -16;
assign rom[82][0] = -19;
assign rom[82][1] = 12;
assign rom[82][2] = 13;
assign rom[82][3] = 20;
assign rom[82][4] = 9;
assign rom[82][5] = -16;
assign rom[82][6] = -11;
assign rom[82][7] = -4;
assign rom[82][8] = -20;
assign rom[82][9] = -20;
assign rom[83][0] = -4;
assign rom[83][1] = -3;
assign rom[83][2] = 3;
assign rom[83][3] = 26;
assign rom[83][4] = -6;
assign rom[83][5] = -15;
assign rom[83][6] = -1;
assign rom[83][7] = -9;
assign rom[83][8] = -19;
assign rom[83][9] = -8;
assign rom[84][0] = -13;
assign rom[84][1] = -10;
assign rom[84][2] = 13;
assign rom[84][3] = 14;
assign rom[84][4] = -6;
assign rom[84][5] = -12;
assign rom[84][6] = 6;
assign rom[84][7] = 0;
assign rom[84][8] = -10;
assign rom[84][9] = -19;
assign rom[85][0] = -5;
assign rom[85][1] = -28;
assign rom[85][2] = 24;
assign rom[85][3] = 17;
assign rom[85][4] = -12;
assign rom[85][5] = -12;
assign rom[85][6] = -3;
assign rom[85][7] = -9;
assign rom[85][8] = -20;
assign rom[85][9] = -25;
assign rom[86][0] = 0;
assign rom[86][1] = -7;
assign rom[86][2] = 24;
assign rom[86][3] = 12;
assign rom[86][4] = -7;
assign rom[86][5] = -20;
assign rom[86][6] = 11;
assign rom[86][7] = -19;
assign rom[86][8] = -11;
assign rom[86][9] = -21;
assign rom[87][0] = -6;
assign rom[87][1] = 3;
assign rom[87][2] = 23;
assign rom[87][3] = 11;
assign rom[87][4] = -18;
assign rom[87][5] = -20;
assign rom[87][6] = -6;
assign rom[87][7] = -10;
assign rom[87][8] = 1;
assign rom[87][9] = -14;
assign rom[88][0] = 5;
assign rom[88][1] = 6;
assign rom[88][2] = 23;
assign rom[88][3] = 16;
assign rom[88][4] = -21;
assign rom[88][5] = -22;
assign rom[88][6] = -3;
assign rom[88][7] = -16;
assign rom[88][8] = 4;
assign rom[88][9] = -10;
assign rom[89][0] = 2;
assign rom[89][1] = 15;
assign rom[89][2] = 26;
assign rom[89][3] = 11;
assign rom[89][4] = -13;
assign rom[89][5] = -12;
assign rom[89][6] = -3;
assign rom[89][7] = -36;
assign rom[89][8] = 10;
assign rom[89][9] = -14;
assign rom[90][0] = 1;
assign rom[90][1] = 17;
assign rom[90][2] = 22;
assign rom[90][3] = -2;
assign rom[90][4] = -21;
assign rom[90][5] = -10;
assign rom[90][6] = -8;
assign rom[90][7] = -33;
assign rom[90][8] = 8;
assign rom[90][9] = -34;
assign rom[91][0] = 13;
assign rom[91][1] = 5;
assign rom[91][2] = 17;
assign rom[91][3] = 6;
assign rom[91][4] = -18;
assign rom[91][5] = -17;
assign rom[91][6] = 5;
assign rom[91][7] = -37;
assign rom[91][8] = 14;
assign rom[91][9] = -43;
assign rom[92][0] = 8;
assign rom[92][1] = -4;
assign rom[92][2] = 30;
assign rom[92][3] = -3;
assign rom[92][4] = -1;
assign rom[92][5] = 0;
assign rom[92][6] = 12;
assign rom[92][7] = -35;
assign rom[92][8] = 7;
assign rom[92][9] = -56;
assign rom[93][0] = 7;
assign rom[93][1] = -16;
assign rom[93][2] = 13;
assign rom[93][3] = 11;
assign rom[93][4] = 16;
assign rom[93][5] = -8;
assign rom[93][6] = 4;
assign rom[93][7] = -41;
assign rom[93][8] = -1;
assign rom[93][9] = -56;
assign rom[94][0] = -4;
assign rom[94][1] = -17;
assign rom[94][2] = 17;
assign rom[94][3] = -8;
assign rom[94][4] = 14;
assign rom[94][5] = 7;
assign rom[94][6] = 17;
assign rom[94][7] = -30;
assign rom[94][8] = 7;
assign rom[94][9] = -42;
assign rom[95][0] = 5;
assign rom[95][1] = 6;
assign rom[95][2] = -2;
assign rom[95][3] = -2;
assign rom[95][4] = 0;
assign rom[95][5] = -2;
assign rom[95][6] = 27;
assign rom[95][7] = -25;
assign rom[95][8] = 6;
assign rom[95][9] = -35;
assign rom[96][0] = -6;
assign rom[96][1] = 2;
assign rom[96][2] = 2;
assign rom[96][3] = -10;
assign rom[96][4] = 2;
assign rom[96][5] = 5;
assign rom[96][6] = 33;
assign rom[96][7] = -27;
assign rom[96][8] = -5;
assign rom[96][9] = -29;
assign rom[97][0] = 1;
assign rom[97][1] = 18;
assign rom[97][2] = -9;
assign rom[97][3] = -21;
assign rom[97][4] = 0;
assign rom[97][5] = 0;
assign rom[97][6] = 17;
assign rom[97][7] = -15;
assign rom[97][8] = -8;
assign rom[97][9] = -31;
assign rom[98][0] = -4;
assign rom[98][1] = 24;
assign rom[98][2] = -18;
assign rom[98][3] = -30;
assign rom[98][4] = 18;
assign rom[98][5] = 10;
assign rom[98][6] = 29;
assign rom[98][7] = -15;
assign rom[98][8] = -12;
assign rom[98][9] = -21;
assign rom[99][0] = -20;
assign rom[99][1] = 8;
assign rom[99][2] = -17;
assign rom[99][3] = -48;
assign rom[99][4] = 12;
assign rom[99][5] = 17;
assign rom[99][6] = 21;
assign rom[99][7] = -9;
assign rom[99][8] = -18;
assign rom[99][9] = -24;
assign rom[100][0] = -24;
assign rom[100][1] = 14;
assign rom[100][2] = -22;
assign rom[100][3] = -28;
assign rom[100][4] = 22;
assign rom[100][5] = 7;
assign rom[100][6] = 30;
assign rom[100][7] = -7;
assign rom[100][8] = -16;
assign rom[100][9] = -25;
assign rom[101][0] = -12;
assign rom[101][1] = 9;
assign rom[101][2] = -12;
assign rom[101][3] = -30;
assign rom[101][4] = 19;
assign rom[101][5] = 16;
assign rom[101][6] = 12;
assign rom[101][7] = 12;
assign rom[101][8] = -18;
assign rom[101][9] = -19;
assign rom[102][0] = -12;
assign rom[102][1] = 7;
assign rom[102][2] = -13;
assign rom[102][3] = -7;
assign rom[102][4] = 12;
assign rom[102][5] = 17;
assign rom[102][6] = 12;
assign rom[102][7] = 13;
assign rom[102][8] = -20;
assign rom[102][9] = -1;
assign rom[103][0] = -7;
assign rom[103][1] = 13;
assign rom[103][2] = 0;
assign rom[103][3] = -15;
assign rom[103][4] = 12;
assign rom[103][5] = 8;
assign rom[103][6] = 4;
assign rom[103][7] = 14;
assign rom[103][8] = -30;
assign rom[103][9] = -5;
assign rom[104][0] = 1;
assign rom[104][1] = 27;
assign rom[104][2] = -4;
assign rom[104][3] = -15;
assign rom[104][4] = -1;
assign rom[104][5] = 7;
assign rom[104][6] = -4;
assign rom[104][7] = 7;
assign rom[104][8] = -26;
assign rom[104][9] = -3;
assign rom[105][0] = -16;
assign rom[105][1] = 21;
assign rom[105][2] = -11;
assign rom[105][3] = 9;
assign rom[105][4] = -2;
assign rom[105][5] = 5;
assign rom[105][6] = -7;
assign rom[105][7] = 17;
assign rom[105][8] = -25;
assign rom[105][9] = -7;
assign rom[106][0] = -4;
assign rom[106][1] = 21;
assign rom[106][2] = -7;
assign rom[106][3] = 18;
assign rom[106][4] = 12;
assign rom[106][5] = -9;
assign rom[106][6] = -14;
assign rom[106][7] = 3;
assign rom[106][8] = -36;
assign rom[106][9] = -6;
assign rom[107][0] = -10;
assign rom[107][1] = 5;
assign rom[107][2] = 12;
assign rom[107][3] = 27;
assign rom[107][4] = 19;
assign rom[107][5] = -27;
assign rom[107][6] = -10;
assign rom[107][7] = 15;
assign rom[107][8] = -21;
assign rom[107][9] = -22;
assign rom[108][0] = -8;
assign rom[108][1] = 2;
assign rom[108][2] = 1;
assign rom[108][3] = 21;
assign rom[108][4] = 1;
assign rom[108][5] = -25;
assign rom[108][6] = -19;
assign rom[108][7] = 1;
assign rom[108][8] = -25;
assign rom[108][9] = -22;
assign rom[109][0] = -10;
assign rom[109][1] = -11;
assign rom[109][2] = 10;
assign rom[109][3] = 26;
assign rom[109][4] = 8;
assign rom[109][5] = -31;
assign rom[109][6] = -14;
assign rom[109][7] = 3;
assign rom[109][8] = -22;
assign rom[109][9] = -32;
assign rom[110][0] = -15;
assign rom[110][1] = -22;
assign rom[110][2] = 12;
assign rom[110][3] = 11;
assign rom[110][4] = -2;
assign rom[110][5] = -19;
assign rom[110][6] = -2;
assign rom[110][7] = -2;
assign rom[110][8] = -16;
assign rom[110][9] = -23;
assign rom[111][0] = -16;
assign rom[111][1] = -23;
assign rom[111][2] = 20;
assign rom[111][3] = 18;
assign rom[111][4] = 12;
assign rom[111][5] = -5;
assign rom[111][6] = -8;
assign rom[111][7] = -7;
assign rom[111][8] = -3;
assign rom[111][9] = -21;
assign rom[112][0] = -9;
assign rom[112][1] = -14;
assign rom[112][2] = 15;
assign rom[112][3] = 18;
assign rom[112][4] = -2;
assign rom[112][5] = 0;
assign rom[112][6] = 2;
assign rom[112][7] = -2;
assign rom[112][8] = -2;
assign rom[112][9] = -19;
assign rom[113][0] = -4;
assign rom[113][1] = -18;
assign rom[113][2] = 17;
assign rom[113][3] = 15;
assign rom[113][4] = -3;
assign rom[113][5] = 6;
assign rom[113][6] = -11;
assign rom[113][7] = -15;
assign rom[113][8] = -4;
assign rom[113][9] = -22;
assign rom[114][0] = 11;
assign rom[114][1] = -3;
assign rom[114][2] = 24;
assign rom[114][3] = 9;
assign rom[114][4] = -12;
assign rom[114][5] = 5;
assign rom[114][6] = -7;
assign rom[114][7] = -15;
assign rom[114][8] = 12;
assign rom[114][9] = -5;
assign rom[115][0] = 3;
assign rom[115][1] = 13;
assign rom[115][2] = 16;
assign rom[115][3] = 5;
assign rom[115][4] = -22;
assign rom[115][5] = -10;
assign rom[115][6] = -11;
assign rom[115][7] = -14;
assign rom[115][8] = 1;
assign rom[115][9] = -20;
assign rom[116][0] = 8;
assign rom[116][1] = 5;
assign rom[116][2] = 19;
assign rom[116][3] = 11;
assign rom[116][4] = -15;
assign rom[116][5] = -7;
assign rom[116][6] = -14;
assign rom[116][7] = -20;
assign rom[116][8] = 19;
assign rom[116][9] = -13;
assign rom[117][0] = 8;
assign rom[117][1] = -10;
assign rom[117][2] = 16;
assign rom[117][3] = 6;
assign rom[117][4] = -13;
assign rom[117][5] = -3;
assign rom[117][6] = -18;
assign rom[117][7] = -19;
assign rom[117][8] = 16;
assign rom[117][9] = -13;
assign rom[118][0] = 16;
assign rom[118][1] = -7;
assign rom[118][2] = 18;
assign rom[118][3] = 9;
assign rom[118][4] = -18;
assign rom[118][5] = -8;
assign rom[118][6] = -4;
assign rom[118][7] = -27;
assign rom[118][8] = 20;
assign rom[118][9] = -16;
assign rom[119][0] = 16;
assign rom[119][1] = -11;
assign rom[119][2] = 14;
assign rom[119][3] = -8;
assign rom[119][4] = 4;
assign rom[119][5] = 6;
assign rom[119][6] = -11;
assign rom[119][7] = -29;
assign rom[119][8] = 14;
assign rom[119][9] = -29;
assign rom[120][0] = 15;
assign rom[120][1] = -17;
assign rom[120][2] = 17;
assign rom[120][3] = -5;
assign rom[120][4] = 7;
assign rom[120][5] = 7;
assign rom[120][6] = -8;
assign rom[120][7] = -17;
assign rom[120][8] = 6;
assign rom[120][9] = -26;
assign rom[121][0] = 18;
assign rom[121][1] = -1;
assign rom[121][2] = -2;
assign rom[121][3] = -7;
assign rom[121][4] = 5;
assign rom[121][5] = 5;
assign rom[121][6] = 7;
assign rom[121][7] = -29;
assign rom[121][8] = 8;
assign rom[121][9] = -16;
assign rom[122][0] = -3;
assign rom[122][1] = -3;
assign rom[122][2] = 8;
assign rom[122][3] = 2;
assign rom[122][4] = -8;
assign rom[122][5] = 9;
assign rom[122][6] = 3;
assign rom[122][7] = -29;
assign rom[122][8] = 3;
assign rom[122][9] = -20;
assign rom[123][0] = 7;
assign rom[123][1] = 15;
assign rom[123][2] = -4;
assign rom[123][3] = -7;
assign rom[123][4] = 2;
assign rom[123][5] = 0;
assign rom[123][6] = 11;
assign rom[123][7] = -12;
assign rom[123][8] = -2;
assign rom[123][9] = -23;
assign rom[124][0] = -1;
assign rom[124][1] = 19;
assign rom[124][2] = -17;
assign rom[124][3] = -33;
assign rom[124][4] = 12;
assign rom[124][5] = 5;
assign rom[124][6] = 0;
assign rom[124][7] = -10;
assign rom[124][8] = -8;
assign rom[124][9] = -30;
assign rom[125][0] = -10;
assign rom[125][1] = 11;
assign rom[125][2] = -32;
assign rom[125][3] = -39;
assign rom[125][4] = 21;
assign rom[125][5] = 10;
assign rom[125][6] = 7;
assign rom[125][7] = -24;
assign rom[125][8] = -15;
assign rom[125][9] = -40;
assign rom[126][0] = -13;
assign rom[126][1] = 6;
assign rom[126][2] = -29;
assign rom[126][3] = -50;
assign rom[126][4] = 34;
assign rom[126][5] = 31;
assign rom[126][6] = 2;
assign rom[126][7] = -19;
assign rom[126][8] = -6;
assign rom[126][9] = -42;
assign rom[127][0] = -15;
assign rom[127][1] = 11;
assign rom[127][2] = -28;
assign rom[127][3] = -40;
assign rom[127][4] = 9;
assign rom[127][5] = 31;
assign rom[127][6] = 4;
assign rom[127][7] = -7;
assign rom[127][8] = -5;
assign rom[127][9] = -20;
assign rom[128][0] = -15;
assign rom[128][1] = 19;
assign rom[128][2] = -11;
assign rom[128][3] = -25;
assign rom[128][4] = -3;
assign rom[128][5] = 31;
assign rom[128][6] = 0;
assign rom[128][7] = 1;
assign rom[128][8] = -5;
assign rom[128][9] = -7;
assign rom[129][0] = -17;
assign rom[129][1] = 22;
assign rom[129][2] = -11;
assign rom[129][3] = -14;
assign rom[129][4] = 11;
assign rom[129][5] = 15;
assign rom[129][6] = -8;
assign rom[129][7] = 4;
assign rom[129][8] = -19;
assign rom[129][9] = -9;
assign rom[130][0] = -13;
assign rom[130][1] = 18;
assign rom[130][2] = 4;
assign rom[130][3] = -4;
assign rom[130][4] = 9;
assign rom[130][5] = 22;
assign rom[130][6] = 0;
assign rom[130][7] = 14;
assign rom[130][8] = -17;
assign rom[130][9] = -13;
assign rom[131][0] = -8;
assign rom[131][1] = 12;
assign rom[131][2] = -8;
assign rom[131][3] = 5;
assign rom[131][4] = 12;
assign rom[131][5] = 13;
assign rom[131][6] = -6;
assign rom[131][7] = 21;
assign rom[131][8] = -30;
assign rom[131][9] = -12;
assign rom[132][0] = -8;
assign rom[132][1] = 22;
assign rom[132][2] = -1;
assign rom[132][3] = 14;
assign rom[132][4] = 10;
assign rom[132][5] = -21;
assign rom[132][6] = -11;
assign rom[132][7] = 17;
assign rom[132][8] = -34;
assign rom[132][9] = -10;
assign rom[133][0] = -16;
assign rom[133][1] = -4;
assign rom[133][2] = 7;
assign rom[133][3] = 28;
assign rom[133][4] = 6;
assign rom[133][5] = -28;
assign rom[133][6] = -12;
assign rom[133][7] = 10;
assign rom[133][8] = -23;
assign rom[133][9] = -24;
assign rom[134][0] = -11;
assign rom[134][1] = -18;
assign rom[134][2] = 11;
assign rom[134][3] = 30;
assign rom[134][4] = 3;
assign rom[134][5] = -17;
assign rom[134][6] = -21;
assign rom[134][7] = 6;
assign rom[134][8] = -18;
assign rom[134][9] = -27;
assign rom[135][0] = -14;
assign rom[135][1] = -16;
assign rom[135][2] = 21;
assign rom[135][3] = 21;
assign rom[135][4] = -1;
assign rom[135][5] = -23;
assign rom[135][6] = -4;
assign rom[135][7] = 7;
assign rom[135][8] = -3;
assign rom[135][9] = -41;
assign rom[136][0] = -13;
assign rom[136][1] = -26;
assign rom[136][2] = 18;
assign rom[136][3] = 9;
assign rom[136][4] = -2;
assign rom[136][5] = 3;
assign rom[136][6] = -8;
assign rom[136][7] = 23;
assign rom[136][8] = -11;
assign rom[136][9] = -35;
assign rom[137][0] = -16;
assign rom[137][1] = -32;
assign rom[137][2] = 9;
assign rom[137][3] = 6;
assign rom[137][4] = 10;
assign rom[137][5] = 7;
assign rom[137][6] = -13;
assign rom[137][7] = 16;
assign rom[137][8] = -2;
assign rom[137][9] = -33;
assign rom[138][0] = -2;
assign rom[138][1] = -20;
assign rom[138][2] = 17;
assign rom[138][3] = 10;
assign rom[138][4] = -3;
assign rom[138][5] = 3;
assign rom[138][6] = -7;
assign rom[138][7] = 25;
assign rom[138][8] = 8;
assign rom[138][9] = -18;
assign rom[139][0] = 5;
assign rom[139][1] = -14;
assign rom[139][2] = -1;
assign rom[139][3] = 12;
assign rom[139][4] = -12;
assign rom[139][5] = 11;
assign rom[139][6] = -12;
assign rom[139][7] = 4;
assign rom[139][8] = 3;
assign rom[139][9] = -10;
assign rom[140][0] = -6;
assign rom[140][1] = -2;
assign rom[140][2] = 10;
assign rom[140][3] = 9;
assign rom[140][4] = -22;
assign rom[140][5] = 8;
assign rom[140][6] = -9;
assign rom[140][7] = -1;
assign rom[140][8] = -6;
assign rom[140][9] = -6;
assign rom[141][0] = -1;
assign rom[141][1] = -12;
assign rom[141][2] = 4;
assign rom[141][3] = 15;
assign rom[141][4] = -13;
assign rom[141][5] = -5;
assign rom[141][6] = -22;
assign rom[141][7] = -2;
assign rom[141][8] = 2;
assign rom[141][9] = 14;
assign rom[142][0] = 4;
assign rom[142][1] = -4;
assign rom[142][2] = 10;
assign rom[142][3] = 9;
assign rom[142][4] = -34;
assign rom[142][5] = 3;
assign rom[142][6] = -20;
assign rom[142][7] = -10;
assign rom[142][8] = 12;
assign rom[142][9] = 21;
assign rom[143][0] = 21;
assign rom[143][1] = -18;
assign rom[143][2] = 4;
assign rom[143][3] = 5;
assign rom[143][4] = -29;
assign rom[143][5] = -6;
assign rom[143][6] = -24;
assign rom[143][7] = -28;
assign rom[143][8] = -2;
assign rom[143][9] = 30;
assign rom[144][0] = 26;
assign rom[144][1] = -17;
assign rom[144][2] = 5;
assign rom[144][3] = 11;
assign rom[144][4] = -35;
assign rom[144][5] = -10;
assign rom[144][6] = -17;
assign rom[144][7] = -24;
assign rom[144][8] = 9;
assign rom[144][9] = 37;
assign rom[145][0] = 14;
assign rom[145][1] = -21;
assign rom[145][2] = 7;
assign rom[145][3] = 1;
assign rom[145][4] = -28;
assign rom[145][5] = -3;
assign rom[145][6] = -13;
assign rom[145][7] = -23;
assign rom[145][8] = 17;
assign rom[145][9] = 34;
assign rom[146][0] = 19;
assign rom[146][1] = -13;
assign rom[146][2] = 10;
assign rom[146][3] = 12;
assign rom[146][4] = -18;
assign rom[146][5] = 10;
assign rom[146][6] = -9;
assign rom[146][7] = -12;
assign rom[146][8] = 10;
assign rom[146][9] = 9;
assign rom[147][0] = 16;
assign rom[147][1] = -2;
assign rom[147][2] = 0;
assign rom[147][3] = 4;
assign rom[147][4] = -22;
assign rom[147][5] = 14;
assign rom[147][6] = -7;
assign rom[147][7] = -19;
assign rom[147][8] = 1;
assign rom[147][9] = 7;
assign rom[148][0] = 12;
assign rom[148][1] = 1;
assign rom[148][2] = -6;
assign rom[148][3] = -3;
assign rom[148][4] = -12;
assign rom[148][5] = 5;
assign rom[148][6] = -11;
assign rom[148][7] = -15;
assign rom[148][8] = -4;
assign rom[148][9] = -13;
assign rom[149][0] = 1;
assign rom[149][1] = 9;
assign rom[149][2] = -1;
assign rom[149][3] = 3;
assign rom[149][4] = -3;
assign rom[149][5] = 15;
assign rom[149][6] = -6;
assign rom[149][7] = -8;
assign rom[149][8] = 7;
assign rom[149][9] = -3;
assign rom[150][0] = 14;
assign rom[150][1] = -2;
assign rom[150][2] = -6;
assign rom[150][3] = -6;
assign rom[150][4] = 10;
assign rom[150][5] = 4;
assign rom[150][6] = -16;
assign rom[150][7] = -4;
assign rom[150][8] = 12;
assign rom[150][9] = -19;
assign rom[151][0] = 8;
assign rom[151][1] = -10;
assign rom[151][2] = -25;
assign rom[151][3] = -25;
assign rom[151][4] = 15;
assign rom[151][5] = 21;
assign rom[151][6] = -7;
assign rom[151][7] = -9;
assign rom[151][8] = 1;
assign rom[151][9] = -31;
assign rom[152][0] = -3;
assign rom[152][1] = -12;
assign rom[152][2] = -30;
assign rom[152][3] = -49;
assign rom[152][4] = 26;
assign rom[152][5] = 26;
assign rom[152][6] = -9;
assign rom[152][7] = -22;
assign rom[152][8] = 5;
assign rom[152][9] = -35;
assign rom[153][0] = -28;
assign rom[153][1] = -14;
assign rom[153][2] = -35;
assign rom[153][3] = -32;
assign rom[153][4] = 21;
assign rom[153][5] = 40;
assign rom[153][6] = -20;
assign rom[153][7] = -14;
assign rom[153][8] = 12;
assign rom[153][9] = -43;
assign rom[154][0] = -32;
assign rom[154][1] = 9;
assign rom[154][2] = -3;
assign rom[154][3] = -18;
assign rom[154][4] = 7;
assign rom[154][5] = 32;
assign rom[154][6] = -4;
assign rom[154][7] = -5;
assign rom[154][8] = -3;
assign rom[154][9] = -20;
assign rom[155][0] = -24;
assign rom[155][1] = 21;
assign rom[155][2] = 0;
assign rom[155][3] = -16;
assign rom[155][4] = 11;
assign rom[155][5] = 20;
assign rom[155][6] = -13;
assign rom[155][7] = -1;
assign rom[155][8] = -14;
assign rom[155][9] = -7;
assign rom[156][0] = -5;
assign rom[156][1] = 15;
assign rom[156][2] = 2;
assign rom[156][3] = -2;
assign rom[156][4] = 6;
assign rom[156][5] = 7;
assign rom[156][6] = -5;
assign rom[156][7] = 24;
assign rom[156][8] = -34;
assign rom[156][9] = -1;
assign rom[157][0] = -13;
assign rom[157][1] = 23;
assign rom[157][2] = 2;
assign rom[157][3] = 9;
assign rom[157][4] = 5;
assign rom[157][5] = -5;
assign rom[157][6] = -16;
assign rom[157][7] = 16;
assign rom[157][8] = -18;
assign rom[157][9] = -14;
assign rom[158][0] = -17;
assign rom[158][1] = 8;
assign rom[158][2] = 14;
assign rom[158][3] = 26;
assign rom[158][4] = -2;
assign rom[158][5] = -35;
assign rom[158][6] = -2;
assign rom[158][7] = 19;
assign rom[158][8] = -27;
assign rom[158][9] = -32;
assign rom[159][0] = -22;
assign rom[159][1] = 6;
assign rom[159][2] = 19;
assign rom[159][3] = 17;
assign rom[159][4] = 8;
assign rom[159][5] = -21;
assign rom[159][6] = -4;
assign rom[159][7] = 15;
assign rom[159][8] = -7;
assign rom[159][9] = -42;
assign rom[160][0] = -12;
assign rom[160][1] = -24;
assign rom[160][2] = 21;
assign rom[160][3] = 29;
assign rom[160][4] = 6;
assign rom[160][5] = -19;
assign rom[160][6] = -5;
assign rom[160][7] = 24;
assign rom[160][8] = -6;
assign rom[160][9] = -34;
assign rom[161][0] = -5;
assign rom[161][1] = -30;
assign rom[161][2] = 19;
assign rom[161][3] = 18;
assign rom[161][4] = 1;
assign rom[161][5] = -14;
assign rom[161][6] = -1;
assign rom[161][7] = 28;
assign rom[161][8] = 6;
assign rom[161][9] = -36;
assign rom[162][0] = -18;
assign rom[162][1] = -27;
assign rom[162][2] = 11;
assign rom[162][3] = 20;
assign rom[162][4] = 0;
assign rom[162][5] = -9;
assign rom[162][6] = -12;
assign rom[162][7] = 26;
assign rom[162][8] = -5;
assign rom[162][9] = -28;
assign rom[163][0] = -9;
assign rom[163][1] = -34;
assign rom[163][2] = 11;
assign rom[163][3] = 18;
assign rom[163][4] = 0;
assign rom[163][5] = 0;
assign rom[163][6] = -4;
assign rom[163][7] = 21;
assign rom[163][8] = -4;
assign rom[163][9] = -19;
assign rom[164][0] = 0;
assign rom[164][1] = -28;
assign rom[164][2] = 3;
assign rom[164][3] = 8;
assign rom[164][4] = -13;
assign rom[164][5] = 1;
assign rom[164][6] = -20;
assign rom[164][7] = 16;
assign rom[164][8] = -1;
assign rom[164][9] = -24;
assign rom[165][0] = -9;
assign rom[165][1] = -25;
assign rom[165][2] = 14;
assign rom[165][3] = 3;
assign rom[165][4] = -17;
assign rom[165][5] = 5;
assign rom[165][6] = -13;
assign rom[165][7] = 28;
assign rom[165][8] = -3;
assign rom[165][9] = -11;
assign rom[166][0] = 7;
assign rom[166][1] = -13;
assign rom[166][2] = 3;
assign rom[166][3] = -2;
assign rom[166][4] = -28;
assign rom[166][5] = 10;
assign rom[166][6] = -20;
assign rom[166][7] = 21;
assign rom[166][8] = -3;
assign rom[166][9] = 1;
assign rom[167][0] = -2;
assign rom[167][1] = -16;
assign rom[167][2] = 14;
assign rom[167][3] = 9;
assign rom[167][4] = -31;
assign rom[167][5] = -2;
assign rom[167][6] = -25;
assign rom[167][7] = 1;
assign rom[167][8] = -2;
assign rom[167][9] = 14;
assign rom[168][0] = 10;
assign rom[168][1] = -4;
assign rom[168][2] = 5;
assign rom[168][3] = 12;
assign rom[168][4] = -31;
assign rom[168][5] = -1;
assign rom[168][6] = -14;
assign rom[168][7] = 6;
assign rom[168][8] = -10;
assign rom[168][9] = 39;
assign rom[169][0] = 2;
assign rom[169][1] = -2;
assign rom[169][2] = 13;
assign rom[169][3] = 7;
assign rom[169][4] = -43;
assign rom[169][5] = -8;
assign rom[169][6] = -8;
assign rom[169][7] = 6;
assign rom[169][8] = -10;
assign rom[169][9] = 38;
assign rom[170][0] = 26;
assign rom[170][1] = -9;
assign rom[170][2] = 1;
assign rom[170][3] = 4;
assign rom[170][4] = -50;
assign rom[170][5] = -9;
assign rom[170][6] = -21;
assign rom[170][7] = -6;
assign rom[170][8] = 7;
assign rom[170][9] = 44;
assign rom[171][0] = 22;
assign rom[171][1] = -15;
assign rom[171][2] = 10;
assign rom[171][3] = 13;
assign rom[171][4] = -43;
assign rom[171][5] = -6;
assign rom[171][6] = -12;
assign rom[171][7] = 10;
assign rom[171][8] = 2;
assign rom[171][9] = 30;
assign rom[172][0] = 24;
assign rom[172][1] = -19;
assign rom[172][2] = -5;
assign rom[172][3] = 10;
assign rom[172][4] = -28;
assign rom[172][5] = -1;
assign rom[172][6] = -31;
assign rom[172][7] = 12;
assign rom[172][8] = 1;
assign rom[172][9] = 14;
assign rom[173][0] = 27;
assign rom[173][1] = -1;
assign rom[173][2] = -2;
assign rom[173][3] = 6;
assign rom[173][4] = -17;
assign rom[173][5] = 3;
assign rom[173][6] = -26;
assign rom[173][7] = 16;
assign rom[173][8] = 14;
assign rom[173][9] = 4;
assign rom[174][0] = 14;
assign rom[174][1] = -5;
assign rom[174][2] = -4;
assign rom[174][3] = 8;
assign rom[174][4] = -5;
assign rom[174][5] = 1;
assign rom[174][6] = -38;
assign rom[174][7] = 16;
assign rom[174][8] = 7;
assign rom[174][9] = 3;
assign rom[175][0] = 15;
assign rom[175][1] = 3;
assign rom[175][2] = -5;
assign rom[175][3] = 4;
assign rom[175][4] = -2;
assign rom[175][5] = 9;
assign rom[175][6] = -21;
assign rom[175][7] = -1;
assign rom[175][8] = 3;
assign rom[175][9] = 2;
assign rom[176][0] = 8;
assign rom[176][1] = -7;
assign rom[176][2] = -2;
assign rom[176][3] = 2;
assign rom[176][4] = -1;
assign rom[176][5] = 8;
assign rom[176][6] = -30;
assign rom[176][7] = 0;
assign rom[176][8] = -1;
assign rom[176][9] = -16;
assign rom[177][0] = 20;
assign rom[177][1] = -19;
assign rom[177][2] = -17;
assign rom[177][3] = -26;
assign rom[177][4] = 20;
assign rom[177][5] = 14;
assign rom[177][6] = -25;
assign rom[177][7] = -9;
assign rom[177][8] = 3;
assign rom[177][9] = -29;
assign rom[178][0] = 6;
assign rom[178][1] = -29;
assign rom[178][2] = -37;
assign rom[178][3] = -49;
assign rom[178][4] = 10;
assign rom[178][5] = 30;
assign rom[178][6] = -29;
assign rom[178][7] = -21;
assign rom[178][8] = 13;
assign rom[178][9] = -33;
assign rom[179][0] = -23;
assign rom[179][1] = -19;
assign rom[179][2] = -40;
assign rom[179][3] = -49;
assign rom[179][4] = 14;
assign rom[179][5] = 53;
assign rom[179][6] = -25;
assign rom[179][7] = -17;
assign rom[179][8] = 2;
assign rom[179][9] = -42;
assign rom[180][0] = -34;
assign rom[180][1] = 3;
assign rom[180][2] = -22;
assign rom[180][3] = -21;
assign rom[180][4] = -2;
assign rom[180][5] = 41;
assign rom[180][6] = -16;
assign rom[180][7] = -17;
assign rom[180][8] = -8;
assign rom[180][9] = -27;
assign rom[181][0] = -19;
assign rom[181][1] = 19;
assign rom[181][2] = -11;
assign rom[181][3] = -17;
assign rom[181][4] = 12;
assign rom[181][5] = 28;
assign rom[181][6] = -1;
assign rom[181][7] = -4;
assign rom[181][8] = -16;
assign rom[181][9] = -9;
assign rom[182][0] = -18;
assign rom[182][1] = 18;
assign rom[182][2] = -12;
assign rom[182][3] = -10;
assign rom[182][4] = 10;
assign rom[182][5] = 9;
assign rom[182][6] = -14;
assign rom[182][7] = 15;
assign rom[182][8] = -25;
assign rom[182][9] = -21;
assign rom[183][0] = -23;
assign rom[183][1] = 18;
assign rom[183][2] = -11;
assign rom[183][3] = 2;
assign rom[183][4] = -11;
assign rom[183][5] = -12;
assign rom[183][6] = -2;
assign rom[183][7] = 34;
assign rom[183][8] = -31;
assign rom[183][9] = -21;
assign rom[184][0] = -26;
assign rom[184][1] = 19;
assign rom[184][2] = 13;
assign rom[184][3] = 12;
assign rom[184][4] = 1;
assign rom[184][5] = -33;
assign rom[184][6] = -18;
assign rom[184][7] = 20;
assign rom[184][8] = -23;
assign rom[184][9] = -36;
assign rom[185][0] = -20;
assign rom[185][1] = 0;
assign rom[185][2] = 8;
assign rom[185][3] = 21;
assign rom[185][4] = -10;
assign rom[185][5] = -33;
assign rom[185][6] = -22;
assign rom[185][7] = 18;
assign rom[185][8] = -2;
assign rom[185][9] = -37;
assign rom[186][0] = -14;
assign rom[186][1] = -16;
assign rom[186][2] = 19;
assign rom[186][3] = 24;
assign rom[186][4] = -8;
assign rom[186][5] = -28;
assign rom[186][6] = -17;
assign rom[186][7] = 15;
assign rom[186][8] = 8;
assign rom[186][9] = -32;
assign rom[187][0] = -9;
assign rom[187][1] = -22;
assign rom[187][2] = 2;
assign rom[187][3] = 7;
assign rom[187][4] = -1;
assign rom[187][5] = -13;
assign rom[187][6] = -15;
assign rom[187][7] = 16;
assign rom[187][8] = -1;
assign rom[187][9] = -29;
assign rom[188][0] = -12;
assign rom[188][1] = -33;
assign rom[188][2] = 2;
assign rom[188][3] = 5;
assign rom[188][4] = -4;
assign rom[188][5] = -6;
assign rom[188][6] = 3;
assign rom[188][7] = 6;
assign rom[188][8] = 15;
assign rom[188][9] = -20;
assign rom[189][0] = -2;
assign rom[189][1] = -36;
assign rom[189][2] = -2;
assign rom[189][3] = -10;
assign rom[189][4] = -15;
assign rom[189][5] = 13;
assign rom[189][6] = -4;
assign rom[189][7] = 17;
assign rom[189][8] = 14;
assign rom[189][9] = -12;
assign rom[190][0] = -13;
assign rom[190][1] = -27;
assign rom[190][2] = 12;
assign rom[190][3] = -1;
assign rom[190][4] = -6;
assign rom[190][5] = 6;
assign rom[190][6] = -22;
assign rom[190][7] = 20;
assign rom[190][8] = 3;
assign rom[190][9] = -5;
assign rom[191][0] = -3;
assign rom[191][1] = -18;
assign rom[191][2] = 11;
assign rom[191][3] = -6;
assign rom[191][4] = -8;
assign rom[191][5] = 14;
assign rom[191][6] = -10;
assign rom[191][7] = 14;
assign rom[191][8] = 10;
assign rom[191][9] = 2;
assign rom[192][0] = 2;
assign rom[192][1] = -11;
assign rom[192][2] = 6;
assign rom[192][3] = -11;
assign rom[192][4] = -10;
assign rom[192][5] = 10;
assign rom[192][6] = -18;
assign rom[192][7] = 11;
assign rom[192][8] = 3;
assign rom[192][9] = 18;
assign rom[193][0] = 6;
assign rom[193][1] = -11;
assign rom[193][2] = 11;
assign rom[193][3] = -21;
assign rom[193][4] = -23;
assign rom[193][5] = -2;
assign rom[193][6] = -10;
assign rom[193][7] = 22;
assign rom[193][8] = 3;
assign rom[193][9] = 10;
assign rom[194][0] = 7;
assign rom[194][1] = -2;
assign rom[194][2] = 6;
assign rom[194][3] = -2;
assign rom[194][4] = -42;
assign rom[194][5] = -3;
assign rom[194][6] = -13;
assign rom[194][7] = 16;
assign rom[194][8] = -1;
assign rom[194][9] = 17;
assign rom[195][0] = 19;
assign rom[195][1] = -1;
assign rom[195][2] = -1;
assign rom[195][3] = 4;
assign rom[195][4] = -45;
assign rom[195][5] = -20;
assign rom[195][6] = -25;
assign rom[195][7] = 19;
assign rom[195][8] = -6;
assign rom[195][9] = 22;
assign rom[196][0] = 17;
assign rom[196][1] = -1;
assign rom[196][2] = 11;
assign rom[196][3] = 24;
assign rom[196][4] = -37;
assign rom[196][5] = -20;
assign rom[196][6] = -15;
assign rom[196][7] = 21;
assign rom[196][8] = -19;
assign rom[196][9] = 12;
assign rom[197][0] = 33;
assign rom[197][1] = 7;
assign rom[197][2] = 10;
assign rom[197][3] = 16;
assign rom[197][4] = -19;
assign rom[197][5] = -11;
assign rom[197][6] = -29;
assign rom[197][7] = 29;
assign rom[197][8] = -11;
assign rom[197][9] = 15;
assign rom[198][0] = 22;
assign rom[198][1] = 2;
assign rom[198][2] = 6;
assign rom[198][3] = 5;
assign rom[198][4] = -8;
assign rom[198][5] = -13;
assign rom[198][6] = -31;
assign rom[198][7] = 26;
assign rom[198][8] = -13;
assign rom[198][9] = 1;
assign rom[199][0] = 25;
assign rom[199][1] = -5;
assign rom[199][2] = -8;
assign rom[199][3] = 11;
assign rom[199][4] = -4;
assign rom[199][5] = -8;
assign rom[199][6] = -38;
assign rom[199][7] = 25;
assign rom[199][8] = 1;
assign rom[199][9] = -9;
assign rom[200][0] = 17;
assign rom[200][1] = -14;
assign rom[200][2] = 5;
assign rom[200][3] = 11;
assign rom[200][4] = -6;
assign rom[200][5] = 6;
assign rom[200][6] = -42;
assign rom[200][7] = 22;
assign rom[200][8] = -2;
assign rom[200][9] = -5;
assign rom[201][0] = 0;
assign rom[201][1] = -12;
assign rom[201][2] = 0;
assign rom[201][3] = 9;
assign rom[201][4] = -12;
assign rom[201][5] = 17;
assign rom[201][6] = -39;
assign rom[201][7] = 17;
assign rom[201][8] = 8;
assign rom[201][9] = -2;
assign rom[202][0] = 7;
assign rom[202][1] = -28;
assign rom[202][2] = 0;
assign rom[202][3] = -1;
assign rom[202][4] = 3;
assign rom[202][5] = 22;
assign rom[202][6] = -29;
assign rom[202][7] = -4;
assign rom[202][8] = 17;
assign rom[202][9] = -22;
assign rom[203][0] = 9;
assign rom[203][1] = -34;
assign rom[203][2] = -23;
assign rom[203][3] = -17;
assign rom[203][4] = 3;
assign rom[203][5] = 27;
assign rom[203][6] = -43;
assign rom[203][7] = -15;
assign rom[203][8] = 4;
assign rom[203][9] = -21;
assign rom[204][0] = 7;
assign rom[204][1] = -38;
assign rom[204][2] = -26;
assign rom[204][3] = -31;
assign rom[204][4] = -5;
assign rom[204][5] = 41;
assign rom[204][6] = -38;
assign rom[204][7] = -14;
assign rom[204][8] = 12;
assign rom[204][9] = -36;
assign rom[205][0] = -15;
assign rom[205][1] = -38;
assign rom[205][2] = -39;
assign rom[205][3] = -41;
assign rom[205][4] = -3;
assign rom[205][5] = 56;
assign rom[205][6] = -31;
assign rom[205][7] = -24;
assign rom[205][8] = 0;
assign rom[205][9] = -44;
assign rom[206][0] = -22;
assign rom[206][1] = -17;
assign rom[206][2] = -15;
assign rom[206][3] = -34;
assign rom[206][4] = -6;
assign rom[206][5] = 60;
assign rom[206][6] = -34;
assign rom[206][7] = -15;
assign rom[206][8] = -13;
assign rom[206][9] = -31;
assign rom[207][0] = -18;
assign rom[207][1] = 18;
assign rom[207][2] = -3;
assign rom[207][3] = -19;
assign rom[207][4] = -4;
assign rom[207][5] = 34;
assign rom[207][6] = -19;
assign rom[207][7] = 8;
assign rom[207][8] = -14;
assign rom[207][9] = -8;
assign rom[208][0] = -11;
assign rom[208][1] = 24;
assign rom[208][2] = -13;
assign rom[208][3] = -6;
assign rom[208][4] = 7;
assign rom[208][5] = 10;
assign rom[208][6] = 4;
assign rom[208][7] = 23;
assign rom[208][8] = -29;
assign rom[208][9] = -24;
assign rom[209][0] = -23;
assign rom[209][1] = 14;
assign rom[209][2] = -9;
assign rom[209][3] = 11;
assign rom[209][4] = -11;
assign rom[209][5] = -12;
assign rom[209][6] = -11;
assign rom[209][7] = 29;
assign rom[209][8] = -28;
assign rom[209][9] = -29;
assign rom[210][0] = -25;
assign rom[210][1] = 3;
assign rom[210][2] = 16;
assign rom[210][3] = 13;
assign rom[210][4] = -16;
assign rom[210][5] = -28;
assign rom[210][6] = -8;
assign rom[210][7] = 31;
assign rom[210][8] = -12;
assign rom[210][9] = -28;
assign rom[211][0] = -11;
assign rom[211][1] = -4;
assign rom[211][2] = 10;
assign rom[211][3] = 19;
assign rom[211][4] = -20;
assign rom[211][5] = -27;
assign rom[211][6] = -6;
assign rom[211][7] = 25;
assign rom[211][8] = -4;
assign rom[211][9] = -19;
assign rom[212][0] = -3;
assign rom[212][1] = -8;
assign rom[212][2] = 7;
assign rom[212][3] = 18;
assign rom[212][4] = -25;
assign rom[212][5] = -12;
assign rom[212][6] = -4;
assign rom[212][7] = 14;
assign rom[212][8] = 10;
assign rom[212][9] = -6;
assign rom[213][0] = -4;
assign rom[213][1] = -20;
assign rom[213][2] = -9;
assign rom[213][3] = 8;
assign rom[213][4] = -15;
assign rom[213][5] = -9;
assign rom[213][6] = -7;
assign rom[213][7] = 3;
assign rom[213][8] = 14;
assign rom[213][9] = -9;
assign rom[214][0] = -1;
assign rom[214][1] = -28;
assign rom[214][2] = -14;
assign rom[214][3] = 0;
assign rom[214][4] = -6;
assign rom[214][5] = 16;
assign rom[214][6] = -7;
assign rom[214][7] = 7;
assign rom[214][8] = 17;
assign rom[214][9] = 6;
assign rom[215][0] = -2;
assign rom[215][1] = -30;
assign rom[215][2] = -8;
assign rom[215][3] = -10;
assign rom[215][4] = -9;
assign rom[215][5] = 20;
assign rom[215][6] = -15;
assign rom[215][7] = 3;
assign rom[215][8] = 12;
assign rom[215][9] = -3;
assign rom[216][0] = 0;
assign rom[216][1] = -11;
assign rom[216][2] = 8;
assign rom[216][3] = -21;
assign rom[216][4] = 5;
assign rom[216][5] = 10;
assign rom[216][6] = -7;
assign rom[216][7] = 6;
assign rom[216][8] = 16;
assign rom[216][9] = 2;
assign rom[217][0] = -9;
assign rom[217][1] = -22;
assign rom[217][2] = -5;
assign rom[217][3] = -29;
assign rom[217][4] = -1;
assign rom[217][5] = 17;
assign rom[217][6] = -12;
assign rom[217][7] = 12;
assign rom[217][8] = 22;
assign rom[217][9] = 8;
assign rom[218][0] = 4;
assign rom[218][1] = -32;
assign rom[218][2] = 3;
assign rom[218][3] = -47;
assign rom[218][4] = 9;
assign rom[218][5] = 19;
assign rom[218][6] = -18;
assign rom[218][7] = 13;
assign rom[218][8] = 17;
assign rom[218][9] = 5;
assign rom[219][0] = -1;
assign rom[219][1] = 5;
assign rom[219][2] = -10;
assign rom[219][3] = -23;
assign rom[219][4] = -3;
assign rom[219][5] = 9;
assign rom[219][6] = -3;
assign rom[219][7] = 10;
assign rom[219][8] = -3;
assign rom[219][9] = 8;
assign rom[220][0] = 14;
assign rom[220][1] = 15;
assign rom[220][2] = -12;
assign rom[220][3] = -9;
assign rom[220][4] = -41;
assign rom[220][5] = -4;
assign rom[220][6] = -7;
assign rom[220][7] = 24;
assign rom[220][8] = -4;
assign rom[220][9] = -13;
assign rom[221][0] = 14;
assign rom[221][1] = 33;
assign rom[221][2] = -2;
assign rom[221][3] = 21;
assign rom[221][4] = -51;
assign rom[221][5] = -17;
assign rom[221][6] = -24;
assign rom[221][7] = 20;
assign rom[221][8] = -23;
assign rom[221][9] = -9;
assign rom[222][0] = -3;
assign rom[222][1] = 31;
assign rom[222][2] = 4;
assign rom[222][3] = 12;
assign rom[222][4] = -32;
assign rom[222][5] = -29;
assign rom[222][6] = -39;
assign rom[222][7] = 40;
assign rom[222][8] = -13;
assign rom[222][9] = -4;
assign rom[223][0] = 8;
assign rom[223][1] = 13;
assign rom[223][2] = 0;
assign rom[223][3] = 25;
assign rom[223][4] = -13;
assign rom[223][5] = -23;
assign rom[223][6] = -33;
assign rom[223][7] = 41;
assign rom[223][8] = -18;
assign rom[223][9] = -12;
assign rom[224][0] = 22;
assign rom[224][1] = 5;
assign rom[224][2] = 0;
assign rom[224][3] = 10;
assign rom[224][4] = -9;
assign rom[224][5] = -16;
assign rom[224][6] = -45;
assign rom[224][7] = 25;
assign rom[224][8] = -1;
assign rom[224][9] = -14;
assign rom[225][0] = 30;
assign rom[225][1] = -16;
assign rom[225][2] = -1;
assign rom[225][3] = 10;
assign rom[225][4] = -6;
assign rom[225][5] = -7;
assign rom[225][6] = -45;
assign rom[225][7] = 18;
assign rom[225][8] = 10;
assign rom[225][9] = -6;
assign rom[226][0] = 22;
assign rom[226][1] = -18;
assign rom[226][2] = 0;
assign rom[226][3] = 21;
assign rom[226][4] = -11;
assign rom[226][5] = -1;
assign rom[226][6] = -36;
assign rom[226][7] = 8;
assign rom[226][8] = -2;
assign rom[226][9] = -7;
assign rom[227][0] = -2;
assign rom[227][1] = -27;
assign rom[227][2] = 5;
assign rom[227][3] = 11;
assign rom[227][4] = -5;
assign rom[227][5] = 2;
assign rom[227][6] = -34;
assign rom[227][7] = 15;
assign rom[227][8] = 12;
assign rom[227][9] = -12;
assign rom[228][0] = 8;
assign rom[228][1] = -41;
assign rom[228][2] = 1;
assign rom[228][3] = 15;
assign rom[228][4] = -9;
assign rom[228][5] = 0;
assign rom[228][6] = -31;
assign rom[228][7] = 12;
assign rom[228][8] = 11;
assign rom[228][9] = -5;
assign rom[229][0] = 13;
assign rom[229][1] = -37;
assign rom[229][2] = -11;
assign rom[229][3] = -13;
assign rom[229][4] = -18;
assign rom[229][5] = 22;
assign rom[229][6] = -21;
assign rom[229][7] = -6;
assign rom[229][8] = 18;
assign rom[229][9] = -16;
assign rom[230][0] = 24;
assign rom[230][1] = -47;
assign rom[230][2] = -17;
assign rom[230][3] = -35;
assign rom[230][4] = -9;
assign rom[230][5] = 48;
assign rom[230][6] = -30;
assign rom[230][7] = -16;
assign rom[230][8] = 15;
assign rom[230][9] = -32;
assign rom[231][0] = -10;
assign rom[231][1] = -36;
assign rom[231][2] = -27;
assign rom[231][3] = -44;
assign rom[231][4] = -17;
assign rom[231][5] = 63;
assign rom[231][6] = -38;
assign rom[231][7] = -30;
assign rom[231][8] = -5;
assign rom[231][9] = -30;
assign rom[232][0] = -32;
assign rom[232][1] = -5;
assign rom[232][2] = -16;
assign rom[232][3] = -32;
assign rom[232][4] = -33;
assign rom[232][5] = 73;
assign rom[232][6] = -20;
assign rom[232][7] = -9;
assign rom[232][8] = -24;
assign rom[232][9] = -20;
assign rom[233][0] = -30;
assign rom[233][1] = 13;
assign rom[233][2] = 3;
assign rom[233][3] = -16;
assign rom[233][4] = -6;
assign rom[233][5] = 60;
assign rom[233][6] = -14;
assign rom[233][7] = 2;
assign rom[233][8] = -22;
assign rom[233][9] = -2;
assign rom[234][0] = -7;
assign rom[234][1] = 27;
assign rom[234][2] = -5;
assign rom[234][3] = -10;
assign rom[234][4] = -8;
assign rom[234][5] = 15;
assign rom[234][6] = -8;
assign rom[234][7] = 37;
assign rom[234][8] = -29;
assign rom[234][9] = -17;
assign rom[235][0] = -19;
assign rom[235][1] = 14;
assign rom[235][2] = -3;
assign rom[235][3] = 11;
assign rom[235][4] = -19;
assign rom[235][5] = 4;
assign rom[235][6] = -14;
assign rom[235][7] = 40;
assign rom[235][8] = -20;
assign rom[235][9] = -27;
assign rom[236][0] = -32;
assign rom[236][1] = 6;
assign rom[236][2] = -2;
assign rom[236][3] = 6;
assign rom[236][4] = -18;
assign rom[236][5] = -12;
assign rom[236][6] = -16;
assign rom[236][7] = 32;
assign rom[236][8] = -2;
assign rom[236][9] = -16;
assign rom[237][0] = -16;
assign rom[237][1] = -1;
assign rom[237][2] = -1;
assign rom[237][3] = 2;
assign rom[237][4] = -10;
assign rom[237][5] = -10;
assign rom[237][6] = -7;
assign rom[237][7] = 25;
assign rom[237][8] = 5;
assign rom[237][9] = -9;
assign rom[238][0] = -12;
assign rom[238][1] = -1;
assign rom[238][2] = -11;
assign rom[238][3] = 2;
assign rom[238][4] = -6;
assign rom[238][5] = 1;
assign rom[238][6] = -7;
assign rom[238][7] = 5;
assign rom[238][8] = 18;
assign rom[238][9] = -1;
assign rom[239][0] = 5;
assign rom[239][1] = -8;
assign rom[239][2] = -29;
assign rom[239][3] = -16;
assign rom[239][4] = -14;
assign rom[239][5] = -5;
assign rom[239][6] = -5;
assign rom[239][7] = 7;
assign rom[239][8] = 25;
assign rom[239][9] = 10;
assign rom[240][0] = -8;
assign rom[240][1] = -15;
assign rom[240][2] = -23;
assign rom[240][3] = -32;
assign rom[240][4] = -4;
assign rom[240][5] = 5;
assign rom[240][6] = 11;
assign rom[240][7] = 3;
assign rom[240][8] = 21;
assign rom[240][9] = 15;
assign rom[241][0] = -11;
assign rom[241][1] = -9;
assign rom[241][2] = -29;
assign rom[241][3] = -28;
assign rom[241][4] = -2;
assign rom[241][5] = 10;
assign rom[241][6] = -7;
assign rom[241][7] = 12;
assign rom[241][8] = 23;
assign rom[241][9] = 6;
assign rom[242][0] = -5;
assign rom[242][1] = -7;
assign rom[242][2] = -29;
assign rom[242][3] = -48;
assign rom[242][4] = 3;
assign rom[242][5] = 11;
assign rom[242][6] = -1;
assign rom[242][7] = 0;
assign rom[242][8] = 18;
assign rom[242][9] = 18;
assign rom[243][0] = 4;
assign rom[243][1] = -26;
assign rom[243][2] = -28;
assign rom[243][3] = -43;
assign rom[243][4] = 8;
assign rom[243][5] = 20;
assign rom[243][6] = 1;
assign rom[243][7] = 7;
assign rom[243][8] = 15;
assign rom[243][9] = 18;
assign rom[244][0] = 6;
assign rom[244][1] = -24;
assign rom[244][2] = -40;
assign rom[244][3] = -39;
assign rom[244][4] = 20;
assign rom[244][5] = 20;
assign rom[244][6] = -5;
assign rom[244][7] = 15;
assign rom[244][8] = 21;
assign rom[244][9] = 10;
assign rom[245][0] = 6;
assign rom[245][1] = -15;
assign rom[245][2] = -39;
assign rom[245][3] = -30;
assign rom[245][4] = -4;
assign rom[245][5] = 30;
assign rom[245][6] = 8;
assign rom[245][7] = 12;
assign rom[245][8] = 15;
assign rom[245][9] = -3;
assign rom[246][0] = -7;
assign rom[246][1] = 15;
assign rom[246][2] = -47;
assign rom[246][3] = -2;
assign rom[246][4] = -30;
assign rom[246][5] = 13;
assign rom[246][6] = -3;
assign rom[246][7] = 21;
assign rom[246][8] = -1;
assign rom[246][9] = -19;
assign rom[247][0] = -17;
assign rom[247][1] = 33;
assign rom[247][2] = -26;
assign rom[247][3] = 7;
assign rom[247][4] = -34;
assign rom[247][5] = -12;
assign rom[247][6] = -31;
assign rom[247][7] = 18;
assign rom[247][8] = -18;
assign rom[247][9] = -18;
assign rom[248][0] = -22;
assign rom[248][1] = 29;
assign rom[248][2] = -5;
assign rom[248][3] = 26;
assign rom[248][4] = -13;
assign rom[248][5] = -12;
assign rom[248][6] = -31;
assign rom[248][7] = 24;
assign rom[248][8] = -18;
assign rom[248][9] = -14;
assign rom[249][0] = -1;
assign rom[249][1] = 18;
assign rom[249][2] = -8;
assign rom[249][3] = 14;
assign rom[249][4] = 8;
assign rom[249][5] = -25;
assign rom[249][6] = -41;
assign rom[249][7] = 35;
assign rom[249][8] = -22;
assign rom[249][9] = -9;
assign rom[250][0] = 4;
assign rom[250][1] = -10;
assign rom[250][2] = -4;
assign rom[250][3] = 19;
assign rom[250][4] = 11;
assign rom[250][5] = -18;
assign rom[250][6] = -39;
assign rom[250][7] = 29;
assign rom[250][8] = 0;
assign rom[250][9] = 0;
assign rom[251][0] = 13;
assign rom[251][1] = -17;
assign rom[251][2] = -8;
assign rom[251][3] = 12;
assign rom[251][4] = -6;
assign rom[251][5] = -23;
assign rom[251][6] = -34;
assign rom[251][7] = 18;
assign rom[251][8] = -2;
assign rom[251][9] = 6;
assign rom[252][0] = 13;
assign rom[252][1] = -13;
assign rom[252][2] = 6;
assign rom[252][3] = 12;
assign rom[252][4] = -2;
assign rom[252][5] = -24;
assign rom[252][6] = -40;
assign rom[252][7] = 15;
assign rom[252][8] = 15;
assign rom[252][9] = 15;
assign rom[253][0] = 4;
assign rom[253][1] = -32;
assign rom[253][2] = -3;
assign rom[253][3] = 15;
assign rom[253][4] = -4;
assign rom[253][5] = -25;
assign rom[253][6] = -19;
assign rom[253][7] = 15;
assign rom[253][8] = 7;
assign rom[253][9] = -1;
assign rom[254][0] = 7;
assign rom[254][1] = -26;
assign rom[254][2] = -14;
assign rom[254][3] = -4;
assign rom[254][4] = -14;
assign rom[254][5] = -28;
assign rom[254][6] = -14;
assign rom[254][7] = -3;
assign rom[254][8] = 14;
assign rom[254][9] = -1;
assign rom[255][0] = 20;
assign rom[255][1] = -45;
assign rom[255][2] = -19;
assign rom[255][3] = -16;
assign rom[255][4] = -26;
assign rom[255][5] = -3;
assign rom[255][6] = -5;
assign rom[255][7] = -11;
assign rom[255][8] = 8;
assign rom[255][9] = -5;
assign rom[256][0] = 35;
assign rom[256][1] = -36;
assign rom[256][2] = -17;
assign rom[256][3] = -24;
assign rom[256][4] = -34;
assign rom[256][5] = 20;
assign rom[256][6] = -7;
assign rom[256][7] = -18;
assign rom[256][8] = 10;
assign rom[256][9] = -22;
assign rom[257][0] = 8;
assign rom[257][1] = -14;
assign rom[257][2] = -12;
assign rom[257][3] = -38;
assign rom[257][4] = -27;
assign rom[257][5] = 64;
assign rom[257][6] = -17;
assign rom[257][7] = -16;
assign rom[257][8] = -4;
assign rom[257][9] = -26;
assign rom[258][0] = -17;
assign rom[258][1] = -2;
assign rom[258][2] = -1;
assign rom[258][3] = -20;
assign rom[258][4] = -34;
assign rom[258][5] = 66;
assign rom[258][6] = -33;
assign rom[258][7] = -12;
assign rom[258][8] = -15;
assign rom[258][9] = -20;
assign rom[259][0] = -24;
assign rom[259][1] = 10;
assign rom[259][2] = -9;
assign rom[259][3] = -10;
assign rom[259][4] = -2;
assign rom[259][5] = 51;
assign rom[259][6] = -14;
assign rom[259][7] = 7;
assign rom[259][8] = -18;
assign rom[259][9] = -2;
assign rom[260][0] = -4;
assign rom[260][1] = 17;
assign rom[260][2] = -9;
assign rom[260][3] = -10;
assign rom[260][4] = -11;
assign rom[260][5] = 13;
assign rom[260][6] = 3;
assign rom[260][7] = 34;
assign rom[260][8] = -17;
assign rom[260][9] = -9;
assign rom[261][0] = -22;
assign rom[261][1] = 11;
assign rom[261][2] = -11;
assign rom[261][3] = -17;
assign rom[261][4] = -7;
assign rom[261][5] = 8;
assign rom[261][6] = 0;
assign rom[261][7] = 35;
assign rom[261][8] = -20;
assign rom[261][9] = -16;
assign rom[262][0] = -24;
assign rom[262][1] = 20;
assign rom[262][2] = -16;
assign rom[262][3] = -3;
assign rom[262][4] = -26;
assign rom[262][5] = 3;
assign rom[262][6] = -4;
assign rom[262][7] = 32;
assign rom[262][8] = -2;
assign rom[262][9] = -1;
assign rom[263][0] = -19;
assign rom[263][1] = -2;
assign rom[263][2] = -31;
assign rom[263][3] = -19;
assign rom[263][4] = -19;
assign rom[263][5] = 6;
assign rom[263][6] = -12;
assign rom[263][7] = 16;
assign rom[263][8] = 7;
assign rom[263][9] = 16;
assign rom[264][0] = -3;
assign rom[264][1] = -8;
assign rom[264][2] = -38;
assign rom[264][3] = -18;
assign rom[264][4] = -2;
assign rom[264][5] = 12;
assign rom[264][6] = 12;
assign rom[264][7] = 5;
assign rom[264][8] = 13;
assign rom[264][9] = 26;
assign rom[265][0] = 5;
assign rom[265][1] = -17;
assign rom[265][2] = -62;
assign rom[265][3] = -45;
assign rom[265][4] = -8;
assign rom[265][5] = 15;
assign rom[265][6] = 15;
assign rom[265][7] = 3;
assign rom[265][8] = 11;
assign rom[265][9] = 12;
assign rom[266][0] = -7;
assign rom[266][1] = -12;
assign rom[266][2] = -58;
assign rom[266][3] = -46;
assign rom[266][4] = 17;
assign rom[266][5] = 8;
assign rom[266][6] = 15;
assign rom[266][7] = 2;
assign rom[266][8] = 29;
assign rom[266][9] = 12;
assign rom[267][0] = -1;
assign rom[267][1] = -12;
assign rom[267][2] = -53;
assign rom[267][3] = -41;
assign rom[267][4] = 11;
assign rom[267][5] = 15;
assign rom[267][6] = 2;
assign rom[267][7] = 0;
assign rom[267][8] = 24;
assign rom[267][9] = 21;
assign rom[268][0] = -3;
assign rom[268][1] = -19;
assign rom[268][2] = -39;
assign rom[268][3] = -25;
assign rom[268][4] = 13;
assign rom[268][5] = 13;
assign rom[268][6] = 3;
assign rom[268][7] = -2;
assign rom[268][8] = 16;
assign rom[268][9] = 18;
assign rom[269][0] = 10;
assign rom[269][1] = -20;
assign rom[269][2] = -49;
assign rom[269][3] = -29;
assign rom[269][4] = 34;
assign rom[269][5] = 14;
assign rom[269][6] = 0;
assign rom[269][7] = 1;
assign rom[269][8] = 1;
assign rom[269][9] = 2;
assign rom[270][0] = 0;
assign rom[270][1] = -36;
assign rom[270][2] = -48;
assign rom[270][3] = -17;
assign rom[270][4] = 34;
assign rom[270][5] = 24;
assign rom[270][6] = 14;
assign rom[270][7] = -1;
assign rom[270][8] = 20;
assign rom[270][9] = -11;
assign rom[271][0] = -10;
assign rom[271][1] = -8;
assign rom[271][2] = -61;
assign rom[271][3] = -9;
assign rom[271][4] = 10;
assign rom[271][5] = 20;
assign rom[271][6] = -2;
assign rom[271][7] = -20;
assign rom[271][8] = 15;
assign rom[271][9] = -4;
assign rom[272][0] = -17;
assign rom[272][1] = 19;
assign rom[272][2] = -58;
assign rom[272][3] = 9;
assign rom[272][4] = -26;
assign rom[272][5] = 16;
assign rom[272][6] = -8;
assign rom[272][7] = -20;
assign rom[272][8] = 10;
assign rom[272][9] = -2;
assign rom[273][0] = -25;
assign rom[273][1] = 51;
assign rom[273][2] = -39;
assign rom[273][3] = 22;
assign rom[273][4] = -25;
assign rom[273][5] = -5;
assign rom[273][6] = -31;
assign rom[273][7] = 0;
assign rom[273][8] = 9;
assign rom[273][9] = 0;
assign rom[274][0] = -43;
assign rom[274][1] = 41;
assign rom[274][2] = -22;
assign rom[274][3] = 14;
assign rom[274][4] = 7;
assign rom[274][5] = -21;
assign rom[274][6] = -24;
assign rom[274][7] = 14;
assign rom[274][8] = -6;
assign rom[274][9] = 13;
assign rom[275][0] = -40;
assign rom[275][1] = 16;
assign rom[275][2] = -14;
assign rom[275][3] = 14;
assign rom[275][4] = 22;
assign rom[275][5] = -26;
assign rom[275][6] = -24;
assign rom[275][7] = 25;
assign rom[275][8] = -14;
assign rom[275][9] = 18;
assign rom[276][0] = -19;
assign rom[276][1] = 2;
assign rom[276][2] = -12;
assign rom[276][3] = 6;
assign rom[276][4] = 16;
assign rom[276][5] = -27;
assign rom[276][6] = -21;
assign rom[276][7] = 27;
assign rom[276][8] = -10;
assign rom[276][9] = 24;
assign rom[277][0] = 6;
assign rom[277][1] = -22;
assign rom[277][2] = 1;
assign rom[277][3] = 6;
assign rom[277][4] = 9;
assign rom[277][5] = -30;
assign rom[277][6] = -17;
assign rom[277][7] = 24;
assign rom[277][8] = -2;
assign rom[277][9] = 15;
assign rom[278][0] = 0;
assign rom[278][1] = -24;
assign rom[278][2] = -2;
assign rom[278][3] = 9;
assign rom[278][4] = -14;
assign rom[278][5] = -46;
assign rom[278][6] = -20;
assign rom[278][7] = 5;
assign rom[278][8] = 7;
assign rom[278][9] = 27;
assign rom[279][0] = 2;
assign rom[279][1] = -23;
assign rom[279][2] = -10;
assign rom[279][3] = -12;
assign rom[279][4] = -9;
assign rom[279][5] = -44;
assign rom[279][6] = -1;
assign rom[279][7] = 1;
assign rom[279][8] = 7;
assign rom[279][9] = 20;
assign rom[280][0] = 16;
assign rom[280][1] = -25;
assign rom[280][2] = -4;
assign rom[280][3] = -13;
assign rom[280][4] = -23;
assign rom[280][5] = -42;
assign rom[280][6] = 13;
assign rom[280][7] = 5;
assign rom[280][8] = 16;
assign rom[280][9] = 21;
assign rom[281][0] = 21;
assign rom[281][1] = -18;
assign rom[281][2] = -25;
assign rom[281][3] = -22;
assign rom[281][4] = -19;
assign rom[281][5] = -43;
assign rom[281][6] = 12;
assign rom[281][7] = -7;
assign rom[281][8] = 27;
assign rom[281][9] = 7;
assign rom[282][0] = 32;
assign rom[282][1] = -17;
assign rom[282][2] = -14;
assign rom[282][3] = -27;
assign rom[282][4] = -22;
assign rom[282][5] = -23;
assign rom[282][6] = 18;
assign rom[282][7] = -16;
assign rom[282][8] = 21;
assign rom[282][9] = -12;
assign rom[283][0] = 10;
assign rom[283][1] = -4;
assign rom[283][2] = -3;
assign rom[283][3] = -21;
assign rom[283][4] = -18;
assign rom[283][5] = 15;
assign rom[283][6] = 9;
assign rom[283][7] = -10;
assign rom[283][8] = 13;
assign rom[283][9] = -22;
assign rom[284][0] = -14;
assign rom[284][1] = 8;
assign rom[284][2] = -1;
assign rom[284][3] = -22;
assign rom[284][4] = -12;
assign rom[284][5] = 52;
assign rom[284][6] = -19;
assign rom[284][7] = -7;
assign rom[284][8] = -3;
assign rom[284][9] = -14;
assign rom[285][0] = -22;
assign rom[285][1] = 14;
assign rom[285][2] = 0;
assign rom[285][3] = -5;
assign rom[285][4] = 7;
assign rom[285][5] = 37;
assign rom[285][6] = -21;
assign rom[285][7] = 15;
assign rom[285][8] = -21;
assign rom[285][9] = -12;
assign rom[286][0] = 0;
assign rom[286][1] = 29;
assign rom[286][2] = -11;
assign rom[286][3] = -11;
assign rom[286][4] = -9;
assign rom[286][5] = 5;
assign rom[286][6] = -11;
assign rom[286][7] = 17;
assign rom[286][8] = -21;
assign rom[286][9] = -4;
assign rom[287][0] = -15;
assign rom[287][1] = 17;
assign rom[287][2] = -14;
assign rom[287][3] = -10;
assign rom[287][4] = -14;
assign rom[287][5] = 2;
assign rom[287][6] = 1;
assign rom[287][7] = 38;
assign rom[287][8] = -17;
assign rom[287][9] = -6;
assign rom[288][0] = -26;
assign rom[288][1] = 24;
assign rom[288][2] = -17;
assign rom[288][3] = -19;
assign rom[288][4] = -13;
assign rom[288][5] = 19;
assign rom[288][6] = -13;
assign rom[288][7] = 26;
assign rom[288][8] = -8;
assign rom[288][9] = -1;
assign rom[289][0] = -10;
assign rom[289][1] = 2;
assign rom[289][2] = -51;
assign rom[289][3] = -24;
assign rom[289][4] = -2;
assign rom[289][5] = 12;
assign rom[289][6] = -11;
assign rom[289][7] = 27;
assign rom[289][8] = 9;
assign rom[289][9] = 15;
assign rom[290][0] = 0;
assign rom[290][1] = -3;
assign rom[290][2] = -65;
assign rom[290][3] = -35;
assign rom[290][4] = -3;
assign rom[290][5] = 0;
assign rom[290][6] = 7;
assign rom[290][7] = 3;
assign rom[290][8] = 12;
assign rom[290][9] = 26;
assign rom[291][0] = 3;
assign rom[291][1] = -13;
assign rom[291][2] = -75;
assign rom[291][3] = -32;
assign rom[291][4] = 12;
assign rom[291][5] = 19;
assign rom[291][6] = 10;
assign rom[291][7] = 0;
assign rom[291][8] = 6;
assign rom[291][9] = 23;
assign rom[292][0] = 3;
assign rom[292][1] = -11;
assign rom[292][2] = -63;
assign rom[292][3] = -37;
assign rom[292][4] = 24;
assign rom[292][5] = 18;
assign rom[292][6] = 6;
assign rom[292][7] = -1;
assign rom[292][8] = 12;
assign rom[292][9] = 8;
assign rom[293][0] = 1;
assign rom[293][1] = 1;
assign rom[293][2] = -51;
assign rom[293][3] = -25;
assign rom[293][4] = 24;
assign rom[293][5] = 11;
assign rom[293][6] = 8;
assign rom[293][7] = -6;
assign rom[293][8] = 10;
assign rom[293][9] = 23;
assign rom[294][0] = -1;
assign rom[294][1] = -27;
assign rom[294][2] = -51;
assign rom[294][3] = -22;
assign rom[294][4] = 25;
assign rom[294][5] = 10;
assign rom[294][6] = 11;
assign rom[294][7] = -10;
assign rom[294][8] = -9;
assign rom[294][9] = 10;
assign rom[295][0] = 4;
assign rom[295][1] = -47;
assign rom[295][2] = -52;
assign rom[295][3] = -12;
assign rom[295][4] = 31;
assign rom[295][5] = 26;
assign rom[295][6] = 11;
assign rom[295][7] = -26;
assign rom[295][8] = 2;
assign rom[295][9] = 1;
assign rom[296][0] = 14;
assign rom[296][1] = -50;
assign rom[296][2] = -45;
assign rom[296][3] = 1;
assign rom[296][4] = 37;
assign rom[296][5] = 27;
assign rom[296][6] = 15;
assign rom[296][7] = -36;
assign rom[296][8] = 4;
assign rom[296][9] = -9;
assign rom[297][0] = 3;
assign rom[297][1] = -9;
assign rom[297][2] = -49;
assign rom[297][3] = -5;
assign rom[297][4] = 20;
assign rom[297][5] = 16;
assign rom[297][6] = 5;
assign rom[297][7] = -58;
assign rom[297][8] = 18;
assign rom[297][9] = 0;
assign rom[298][0] = -23;
assign rom[298][1] = 36;
assign rom[298][2] = -41;
assign rom[298][3] = 15;
assign rom[298][4] = -10;
assign rom[298][5] = 18;
assign rom[298][6] = -18;
assign rom[298][7] = -45;
assign rom[298][8] = 16;
assign rom[298][9] = 12;
assign rom[299][0] = -47;
assign rom[299][1] = 45;
assign rom[299][2] = -37;
assign rom[299][3] = 7;
assign rom[299][4] = -13;
assign rom[299][5] = 4;
assign rom[299][6] = -15;
assign rom[299][7] = -40;
assign rom[299][8] = 9;
assign rom[299][9] = 14;
assign rom[300][0] = -50;
assign rom[300][1] = 30;
assign rom[300][2] = -28;
assign rom[300][3] = 8;
assign rom[300][4] = 20;
assign rom[300][5] = -22;
assign rom[300][6] = -11;
assign rom[300][7] = 4;
assign rom[300][8] = 13;
assign rom[300][9] = 16;
assign rom[301][0] = -35;
assign rom[301][1] = 12;
assign rom[301][2] = -19;
assign rom[301][3] = 20;
assign rom[301][4] = 24;
assign rom[301][5] = -19;
assign rom[301][6] = -3;
assign rom[301][7] = 8;
assign rom[301][8] = -1;
assign rom[301][9] = 19;
assign rom[302][0] = -27;
assign rom[302][1] = -18;
assign rom[302][2] = -22;
assign rom[302][3] = 15;
assign rom[302][4] = 15;
assign rom[302][5] = -30;
assign rom[302][6] = -7;
assign rom[302][7] = 19;
assign rom[302][8] = 1;
assign rom[302][9] = 19;
assign rom[303][0] = -12;
assign rom[303][1] = -14;
assign rom[303][2] = -7;
assign rom[303][3] = -4;
assign rom[303][4] = -1;
assign rom[303][5] = -30;
assign rom[303][6] = -13;
assign rom[303][7] = 8;
assign rom[303][8] = -5;
assign rom[303][9] = 35;
assign rom[304][0] = -13;
assign rom[304][1] = -14;
assign rom[304][2] = -3;
assign rom[304][3] = -3;
assign rom[304][4] = 4;
assign rom[304][5] = -26;
assign rom[304][6] = -5;
assign rom[304][7] = 1;
assign rom[304][8] = -3;
assign rom[304][9] = 24;
assign rom[305][0] = -7;
assign rom[305][1] = -21;
assign rom[305][2] = 1;
assign rom[305][3] = -33;
assign rom[305][4] = -7;
assign rom[305][5] = -33;
assign rom[305][6] = 3;
assign rom[305][7] = 4;
assign rom[305][8] = 17;
assign rom[305][9] = 22;
assign rom[306][0] = 5;
assign rom[306][1] = -5;
assign rom[306][2] = -21;
assign rom[306][3] = -41;
assign rom[306][4] = -6;
assign rom[306][5] = -53;
assign rom[306][6] = 11;
assign rom[306][7] = -11;
assign rom[306][8] = 16;
assign rom[306][9] = 17;
assign rom[307][0] = 28;
assign rom[307][1] = -15;
assign rom[307][2] = -35;
assign rom[307][3] = -44;
assign rom[307][4] = -3;
assign rom[307][5] = -67;
assign rom[307][6] = 34;
assign rom[307][7] = 0;
assign rom[307][8] = 10;
assign rom[307][9] = 5;
assign rom[308][0] = 29;
assign rom[308][1] = -2;
assign rom[308][2] = -23;
assign rom[308][3] = -42;
assign rom[308][4] = -19;
assign rom[308][5] = -56;
assign rom[308][6] = 29;
assign rom[308][7] = -5;
assign rom[308][8] = 24;
assign rom[308][9] = -9;
assign rom[309][0] = 10;
assign rom[309][1] = 19;
assign rom[309][2] = -5;
assign rom[309][3] = -14;
assign rom[309][4] = -13;
assign rom[309][5] = -41;
assign rom[309][6] = 11;
assign rom[309][7] = -2;
assign rom[309][8] = 27;
assign rom[309][9] = -19;
assign rom[310][0] = -1;
assign rom[310][1] = 21;
assign rom[310][2] = 10;
assign rom[310][3] = -23;
assign rom[310][4] = 7;
assign rom[310][5] = 7;
assign rom[310][6] = -16;
assign rom[310][7] = -3;
assign rom[310][8] = 7;
assign rom[310][9] = -12;
assign rom[311][0] = -13;
assign rom[311][1] = 16;
assign rom[311][2] = 5;
assign rom[311][3] = -21;
assign rom[311][4] = 2;
assign rom[311][5] = 25;
assign rom[311][6] = -23;
assign rom[311][7] = 8;
assign rom[311][8] = -13;
assign rom[311][9] = -2;
assign rom[312][0] = -4;
assign rom[312][1] = 29;
assign rom[312][2] = -15;
assign rom[312][3] = -7;
assign rom[312][4] = 1;
assign rom[312][5] = 17;
assign rom[312][6] = 3;
assign rom[312][7] = 21;
assign rom[312][8] = -24;
assign rom[312][9] = -3;
assign rom[313][0] = -9;
assign rom[313][1] = 12;
assign rom[313][2] = -4;
assign rom[313][3] = 0;
assign rom[313][4] = -6;
assign rom[313][5] = 13;
assign rom[313][6] = -10;
assign rom[313][7] = 21;
assign rom[313][8] = -25;
assign rom[313][9] = -1;
assign rom[314][0] = -22;
assign rom[314][1] = 11;
assign rom[314][2] = -32;
assign rom[314][3] = -17;
assign rom[314][4] = 3;
assign rom[314][5] = 18;
assign rom[314][6] = -15;
assign rom[314][7] = 33;
assign rom[314][8] = -21;
assign rom[314][9] = 12;
assign rom[315][0] = 3;
assign rom[315][1] = 2;
assign rom[315][2] = -50;
assign rom[315][3] = -20;
assign rom[315][4] = 11;
assign rom[315][5] = 6;
assign rom[315][6] = -11;
assign rom[315][7] = 17;
assign rom[315][8] = -13;
assign rom[315][9] = 19;
assign rom[316][0] = 0;
assign rom[316][1] = 6;
assign rom[316][2] = -55;
assign rom[316][3] = -33;
assign rom[316][4] = 18;
assign rom[316][5] = -8;
assign rom[316][6] = 19;
assign rom[316][7] = 10;
assign rom[316][8] = -9;
assign rom[316][9] = 24;
assign rom[317][0] = 17;
assign rom[317][1] = -11;
assign rom[317][2] = -48;
assign rom[317][3] = -25;
assign rom[317][4] = 17;
assign rom[317][5] = -5;
assign rom[317][6] = 13;
assign rom[317][7] = 4;
assign rom[317][8] = -9;
assign rom[317][9] = 12;
assign rom[318][0] = 14;
assign rom[318][1] = -3;
assign rom[318][2] = -40;
assign rom[318][3] = -22;
assign rom[318][4] = 19;
assign rom[318][5] = 2;
assign rom[318][6] = 3;
assign rom[318][7] = -5;
assign rom[318][8] = -9;
assign rom[318][9] = 6;
assign rom[319][0] = 4;
assign rom[319][1] = -13;
assign rom[319][2] = -37;
assign rom[319][3] = -20;
assign rom[319][4] = 22;
assign rom[319][5] = 19;
assign rom[319][6] = 12;
assign rom[319][7] = 1;
assign rom[319][8] = -13;
assign rom[319][9] = 15;
assign rom[320][0] = 14;
assign rom[320][1] = -31;
assign rom[320][2] = -26;
assign rom[320][3] = -5;
assign rom[320][4] = 28;
assign rom[320][5] = 8;
assign rom[320][6] = 17;
assign rom[320][7] = -16;
assign rom[320][8] = -16;
assign rom[320][9] = 0;
assign rom[321][0] = 18;
assign rom[321][1] = -37;
assign rom[321][2] = -22;
assign rom[321][3] = -12;
assign rom[321][4] = 34;
assign rom[321][5] = 22;
assign rom[321][6] = 14;
assign rom[321][7] = -39;
assign rom[321][8] = -13;
assign rom[321][9] = -8;
assign rom[322][0] = 10;
assign rom[322][1] = -41;
assign rom[322][2] = -17;
assign rom[322][3] = 9;
assign rom[322][4] = 34;
assign rom[322][5] = 21;
assign rom[322][6] = 14;
assign rom[322][7] = -58;
assign rom[322][8] = 1;
assign rom[322][9] = 4;
assign rom[323][0] = -2;
assign rom[323][1] = 1;
assign rom[323][2] = -20;
assign rom[323][3] = 10;
assign rom[323][4] = 27;
assign rom[323][5] = 13;
assign rom[323][6] = 0;
assign rom[323][7] = -73;
assign rom[323][8] = 14;
assign rom[323][9] = -6;
assign rom[324][0] = -37;
assign rom[324][1] = 36;
assign rom[324][2] = -11;
assign rom[324][3] = 1;
assign rom[324][4] = -9;
assign rom[324][5] = 4;
assign rom[324][6] = -5;
assign rom[324][7] = -65;
assign rom[324][8] = 29;
assign rom[324][9] = 12;
assign rom[325][0] = -60;
assign rom[325][1] = 31;
assign rom[325][2] = -25;
assign rom[325][3] = 13;
assign rom[325][4] = -10;
assign rom[325][5] = -6;
assign rom[325][6] = 4;
assign rom[325][7] = -28;
assign rom[325][8] = 18;
assign rom[325][9] = 20;
assign rom[326][0] = -65;
assign rom[326][1] = 26;
assign rom[326][2] = -22;
assign rom[326][3] = -2;
assign rom[326][4] = 9;
assign rom[326][5] = -34;
assign rom[326][6] = 7;
assign rom[326][7] = -15;
assign rom[326][8] = 13;
assign rom[326][9] = 26;
assign rom[327][0] = -45;
assign rom[327][1] = 5;
assign rom[327][2] = -22;
assign rom[327][3] = 2;
assign rom[327][4] = 29;
assign rom[327][5] = -26;
assign rom[327][6] = -2;
assign rom[327][7] = 16;
assign rom[327][8] = 8;
assign rom[327][9] = 30;
assign rom[328][0] = -33;
assign rom[328][1] = -22;
assign rom[328][2] = -7;
assign rom[328][3] = 2;
assign rom[328][4] = 22;
assign rom[328][5] = -15;
assign rom[328][6] = 3;
assign rom[328][7] = 14;
assign rom[328][8] = 0;
assign rom[328][9] = 31;
assign rom[329][0] = -12;
assign rom[329][1] = -24;
assign rom[329][2] = -9;
assign rom[329][3] = 3;
assign rom[329][4] = 20;
assign rom[329][5] = -20;
assign rom[329][6] = -16;
assign rom[329][7] = 7;
assign rom[329][8] = -5;
assign rom[329][9] = 29;
assign rom[330][0] = -2;
assign rom[330][1] = -31;
assign rom[330][2] = -12;
assign rom[330][3] = -12;
assign rom[330][4] = 9;
assign rom[330][5] = -5;
assign rom[330][6] = -2;
assign rom[330][7] = 5;
assign rom[330][8] = -3;
assign rom[330][9] = 24;
assign rom[331][0] = -15;
assign rom[331][1] = -26;
assign rom[331][2] = -3;
assign rom[331][3] = -16;
assign rom[331][4] = 19;
assign rom[331][5] = -14;
assign rom[331][6] = -5;
assign rom[331][7] = 6;
assign rom[331][8] = -12;
assign rom[331][9] = 9;
assign rom[332][0] = 7;
assign rom[332][1] = -6;
assign rom[332][2] = -27;
assign rom[332][3] = -23;
assign rom[332][4] = 4;
assign rom[332][5] = -14;
assign rom[332][6] = 25;
assign rom[332][7] = -4;
assign rom[332][8] = -12;
assign rom[332][9] = 7;
assign rom[333][0] = 24;
assign rom[333][1] = -8;
assign rom[333][2] = -32;
assign rom[333][3] = -39;
assign rom[333][4] = 2;
assign rom[333][5] = -42;
assign rom[333][6] = 24;
assign rom[333][7] = 6;
assign rom[333][8] = -7;
assign rom[333][9] = -4;
assign rom[334][0] = 30;
assign rom[334][1] = 2;
assign rom[334][2] = -17;
assign rom[334][3] = -27;
assign rom[334][4] = -10;
assign rom[334][5] = -51;
assign rom[334][6] = 31;
assign rom[334][7] = 2;
assign rom[334][8] = 0;
assign rom[334][9] = -28;
assign rom[335][0] = 26;
assign rom[335][1] = 12;
assign rom[335][2] = -1;
assign rom[335][3] = -19;
assign rom[335][4] = 5;
assign rom[335][5] = -36;
assign rom[335][6] = 23;
assign rom[335][7] = 4;
assign rom[335][8] = 2;
assign rom[335][9] = -29;
assign rom[336][0] = 12;
assign rom[336][1] = 20;
assign rom[336][2] = 3;
assign rom[336][3] = -11;
assign rom[336][4] = 2;
assign rom[336][5] = -11;
assign rom[336][6] = -3;
assign rom[336][7] = 9;
assign rom[336][8] = -11;
assign rom[336][9] = -8;
assign rom[337][0] = -6;
assign rom[337][1] = 24;
assign rom[337][2] = 11;
assign rom[337][3] = -12;
assign rom[337][4] = 13;
assign rom[337][5] = 8;
assign rom[337][6] = -20;
assign rom[337][7] = 10;
assign rom[337][8] = -15;
assign rom[337][9] = -3;
assign rom[338][0] = -3;
assign rom[338][1] = 22;
assign rom[338][2] = -4;
assign rom[338][3] = -12;
assign rom[338][4] = 11;
assign rom[338][5] = 20;
assign rom[338][6] = -1;
assign rom[338][7] = 13;
assign rom[338][8] = -23;
assign rom[338][9] = -13;
assign rom[339][0] = -16;
assign rom[339][1] = 29;
assign rom[339][2] = -5;
assign rom[339][3] = -12;
assign rom[339][4] = 9;
assign rom[339][5] = 3;
assign rom[339][6] = 0;
assign rom[339][7] = 11;
assign rom[339][8] = -15;
assign rom[339][9] = -3;
assign rom[340][0] = -10;
assign rom[340][1] = 17;
assign rom[340][2] = -16;
assign rom[340][3] = 4;
assign rom[340][4] = 2;
assign rom[340][5] = 11;
assign rom[340][6] = -32;
assign rom[340][7] = 8;
assign rom[340][8] = -29;
assign rom[340][9] = 15;
assign rom[341][0] = -1;
assign rom[341][1] = 12;
assign rom[341][2] = -15;
assign rom[341][3] = -5;
assign rom[341][4] = 19;
assign rom[341][5] = -17;
assign rom[341][6] = -4;
assign rom[341][7] = -2;
assign rom[341][8] = -30;
assign rom[341][9] = 12;
assign rom[342][0] = 16;
assign rom[342][1] = -11;
assign rom[342][2] = -36;
assign rom[342][3] = -21;
assign rom[342][4] = 28;
assign rom[342][5] = -14;
assign rom[342][6] = 13;
assign rom[342][7] = 2;
assign rom[342][8] = -13;
assign rom[342][9] = 12;
assign rom[343][0] = 10;
assign rom[343][1] = -4;
assign rom[343][2] = -30;
assign rom[343][3] = -23;
assign rom[343][4] = 22;
assign rom[343][5] = -12;
assign rom[343][6] = 4;
assign rom[343][7] = -3;
assign rom[343][8] = -20;
assign rom[343][9] = 17;
assign rom[344][0] = 15;
assign rom[344][1] = -4;
assign rom[344][2] = -22;
assign rom[344][3] = -20;
assign rom[344][4] = 31;
assign rom[344][5] = -11;
assign rom[344][6] = 10;
assign rom[344][7] = -3;
assign rom[344][8] = -25;
assign rom[344][9] = -4;
assign rom[345][0] = 15;
assign rom[345][1] = -17;
assign rom[345][2] = -15;
assign rom[345][3] = -18;
assign rom[345][4] = 24;
assign rom[345][5] = 15;
assign rom[345][6] = 6;
assign rom[345][7] = -19;
assign rom[345][8] = -30;
assign rom[345][9] = 8;
assign rom[346][0] = 7;
assign rom[346][1] = -25;
assign rom[346][2] = 5;
assign rom[346][3] = -9;
assign rom[346][4] = 25;
assign rom[346][5] = 6;
assign rom[346][6] = 17;
assign rom[346][7] = -26;
assign rom[346][8] = -22;
assign rom[346][9] = -6;
assign rom[347][0] = 6;
assign rom[347][1] = -44;
assign rom[347][2] = 11;
assign rom[347][3] = 3;
assign rom[347][4] = 35;
assign rom[347][5] = 20;
assign rom[347][6] = 15;
assign rom[347][7] = -37;
assign rom[347][8] = -15;
assign rom[347][9] = 1;
assign rom[348][0] = -3;
assign rom[348][1] = -31;
assign rom[348][2] = 12;
assign rom[348][3] = -5;
assign rom[348][4] = 31;
assign rom[348][5] = 11;
assign rom[348][6] = 17;
assign rom[348][7] = -51;
assign rom[348][8] = 14;
assign rom[348][9] = -1;
assign rom[349][0] = -13;
assign rom[349][1] = 12;
assign rom[349][2] = 4;
assign rom[349][3] = 9;
assign rom[349][4] = 18;
assign rom[349][5] = 12;
assign rom[349][6] = -1;
assign rom[349][7] = -66;
assign rom[349][8] = 19;
assign rom[349][9] = 0;
assign rom[350][0] = -48;
assign rom[350][1] = 37;
assign rom[350][2] = 0;
assign rom[350][3] = 3;
assign rom[350][4] = -3;
assign rom[350][5] = -5;
assign rom[350][6] = 7;
assign rom[350][7] = -46;
assign rom[350][8] = 30;
assign rom[350][9] = -5;
assign rom[351][0] = -59;
assign rom[351][1] = 45;
assign rom[351][2] = -4;
assign rom[351][3] = 8;
assign rom[351][4] = 11;
assign rom[351][5] = -17;
assign rom[351][6] = 14;
assign rom[351][7] = -28;
assign rom[351][8] = 7;
assign rom[351][9] = 2;
assign rom[352][0] = -54;
assign rom[352][1] = 15;
assign rom[352][2] = -7;
assign rom[352][3] = 3;
assign rom[352][4] = 27;
assign rom[352][5] = -24;
assign rom[352][6] = 9;
assign rom[352][7] = 2;
assign rom[352][8] = 18;
assign rom[352][9] = 17;
assign rom[353][0] = -43;
assign rom[353][1] = -9;
assign rom[353][2] = -1;
assign rom[353][3] = 1;
assign rom[353][4] = 35;
assign rom[353][5] = -21;
assign rom[353][6] = 4;
assign rom[353][7] = 15;
assign rom[353][8] = -4;
assign rom[353][9] = 23;
assign rom[354][0] = -13;
assign rom[354][1] = -19;
assign rom[354][2] = -9;
assign rom[354][3] = -6;
assign rom[354][4] = 19;
assign rom[354][5] = -23;
assign rom[354][6] = -14;
assign rom[354][7] = 7;
assign rom[354][8] = -3;
assign rom[354][9] = 26;
assign rom[355][0] = -7;
assign rom[355][1] = -28;
assign rom[355][2] = -10;
assign rom[355][3] = 2;
assign rom[355][4] = 26;
assign rom[355][5] = -2;
assign rom[355][6] = -18;
assign rom[355][7] = 17;
assign rom[355][8] = -6;
assign rom[355][9] = 12;
assign rom[356][0] = -7;
assign rom[356][1] = -29;
assign rom[356][2] = -18;
assign rom[356][3] = -5;
assign rom[356][4] = 12;
assign rom[356][5] = 1;
assign rom[356][6] = 1;
assign rom[356][7] = 29;
assign rom[356][8] = -22;
assign rom[356][9] = -1;
assign rom[357][0] = 4;
assign rom[357][1] = -24;
assign rom[357][2] = -15;
assign rom[357][3] = -1;
assign rom[357][4] = 17;
assign rom[357][5] = -9;
assign rom[357][6] = 7;
assign rom[357][7] = 12;
assign rom[357][8] = -28;
assign rom[357][9] = -11;
assign rom[358][0] = 9;
assign rom[358][1] = -11;
assign rom[358][2] = -24;
assign rom[358][3] = -18;
assign rom[358][4] = 6;
assign rom[358][5] = -13;
assign rom[358][6] = 20;
assign rom[358][7] = 16;
assign rom[358][8] = -16;
assign rom[358][9] = -20;
assign rom[359][0] = 27;
assign rom[359][1] = -2;
assign rom[359][2] = -20;
assign rom[359][3] = -6;
assign rom[359][4] = 13;
assign rom[359][5] = -14;
assign rom[359][6] = 30;
assign rom[359][7] = 8;
assign rom[359][8] = -17;
assign rom[359][9] = -30;
assign rom[360][0] = 23;
assign rom[360][1] = -4;
assign rom[360][2] = -8;
assign rom[360][3] = -10;
assign rom[360][4] = 8;
assign rom[360][5] = -27;
assign rom[360][6] = 30;
assign rom[360][7] = -6;
assign rom[360][8] = -12;
assign rom[360][9] = -35;
assign rom[361][0] = 24;
assign rom[361][1] = 10;
assign rom[361][2] = 9;
assign rom[361][3] = -8;
assign rom[361][4] = -7;
assign rom[361][5] = -17;
assign rom[361][6] = 17;
assign rom[361][7] = 0;
assign rom[361][8] = -19;
assign rom[361][9] = -30;
assign rom[362][0] = 6;
assign rom[362][1] = 22;
assign rom[362][2] = 26;
assign rom[362][3] = -14;
assign rom[362][4] = 1;
assign rom[362][5] = 1;
assign rom[362][6] = -8;
assign rom[362][7] = 14;
assign rom[362][8] = -24;
assign rom[362][9] = -16;
assign rom[363][0] = -3;
assign rom[363][1] = 26;
assign rom[363][2] = 13;
assign rom[363][3] = -21;
assign rom[363][4] = 4;
assign rom[363][5] = 16;
assign rom[363][6] = -10;
assign rom[363][7] = 5;
assign rom[363][8] = -28;
assign rom[363][9] = -13;
assign rom[364][0] = -2;
assign rom[364][1] = 14;
assign rom[364][2] = -4;
assign rom[364][3] = -3;
assign rom[364][4] = 14;
assign rom[364][5] = 8;
assign rom[364][6] = 6;
assign rom[364][7] = 15;
assign rom[364][8] = -16;
assign rom[364][9] = -1;
assign rom[365][0] = -17;
assign rom[365][1] = 17;
assign rom[365][2] = -4;
assign rom[365][3] = 11;
assign rom[365][4] = 7;
assign rom[365][5] = 12;
assign rom[365][6] = -9;
assign rom[365][7] = 17;
assign rom[365][8] = -32;
assign rom[365][9] = 0;
assign rom[366][0] = -7;
assign rom[366][1] = 11;
assign rom[366][2] = 2;
assign rom[366][3] = 4;
assign rom[366][4] = -6;
assign rom[366][5] = 7;
assign rom[366][6] = -36;
assign rom[366][7] = 3;
assign rom[366][8] = -38;
assign rom[366][9] = 9;
assign rom[367][0] = 17;
assign rom[367][1] = 1;
assign rom[367][2] = -4;
assign rom[367][3] = -10;
assign rom[367][4] = 14;
assign rom[367][5] = -18;
assign rom[367][6] = -25;
assign rom[367][7] = -10;
assign rom[367][8] = -31;
assign rom[367][9] = 9;
assign rom[368][0] = 15;
assign rom[368][1] = -13;
assign rom[368][2] = 4;
assign rom[368][3] = -19;
assign rom[368][4] = 13;
assign rom[368][5] = -33;
assign rom[368][6] = -3;
assign rom[368][7] = 1;
assign rom[368][8] = -32;
assign rom[368][9] = -4;
assign rom[369][0] = 5;
assign rom[369][1] = -21;
assign rom[369][2] = 7;
assign rom[369][3] = -19;
assign rom[369][4] = 18;
assign rom[369][5] = -22;
assign rom[369][6] = 2;
assign rom[369][7] = -16;
assign rom[369][8] = -20;
assign rom[369][9] = 9;
assign rom[370][0] = 17;
assign rom[370][1] = -11;
assign rom[370][2] = 6;
assign rom[370][3] = -32;
assign rom[370][4] = 29;
assign rom[370][5] = -15;
assign rom[370][6] = 10;
assign rom[370][7] = -16;
assign rom[370][8] = -21;
assign rom[370][9] = 5;
assign rom[371][0] = 14;
assign rom[371][1] = -12;
assign rom[371][2] = -3;
assign rom[371][3] = -31;
assign rom[371][4] = 31;
assign rom[371][5] = -9;
assign rom[371][6] = 12;
assign rom[371][7] = -27;
assign rom[371][8] = -18;
assign rom[371][9] = 7;
assign rom[372][0] = 18;
assign rom[372][1] = -31;
assign rom[372][2] = 8;
assign rom[372][3] = -20;
assign rom[372][4] = 12;
assign rom[372][5] = 3;
assign rom[372][6] = 20;
assign rom[372][7] = -33;
assign rom[372][8] = -7;
assign rom[372][9] = 8;
assign rom[373][0] = 19;
assign rom[373][1] = -28;
assign rom[373][2] = 14;
assign rom[373][3] = -6;
assign rom[373][4] = 18;
assign rom[373][5] = 9;
assign rom[373][6] = 23;
assign rom[373][7] = -29;
assign rom[373][8] = -6;
assign rom[373][9] = 7;
assign rom[374][0] = -13;
assign rom[374][1] = -10;
assign rom[374][2] = 9;
assign rom[374][3] = 0;
assign rom[374][4] = 12;
assign rom[374][5] = 7;
assign rom[374][6] = 12;
assign rom[374][7] = -45;
assign rom[374][8] = 21;
assign rom[374][9] = 0;
assign rom[375][0] = -24;
assign rom[375][1] = 8;
assign rom[375][2] = 23;
assign rom[375][3] = 5;
assign rom[375][4] = 0;
assign rom[375][5] = -10;
assign rom[375][6] = 5;
assign rom[375][7] = -53;
assign rom[375][8] = 15;
assign rom[375][9] = -18;
assign rom[376][0] = -43;
assign rom[376][1] = 40;
assign rom[376][2] = 11;
assign rom[376][3] = 3;
assign rom[376][4] = 14;
assign rom[376][5] = -20;
assign rom[376][6] = 15;
assign rom[376][7] = -36;
assign rom[376][8] = 25;
assign rom[376][9] = -12;
assign rom[377][0] = -68;
assign rom[377][1] = 32;
assign rom[377][2] = 1;
assign rom[377][3] = -6;
assign rom[377][4] = 29;
assign rom[377][5] = -26;
assign rom[377][6] = 2;
assign rom[377][7] = 0;
assign rom[377][8] = 14;
assign rom[377][9] = 3;
assign rom[378][0] = -49;
assign rom[378][1] = 14;
assign rom[378][2] = -5;
assign rom[378][3] = -14;
assign rom[378][4] = 25;
assign rom[378][5] = -17;
assign rom[378][6] = 4;
assign rom[378][7] = 0;
assign rom[378][8] = 1;
assign rom[378][9] = 4;
assign rom[379][0] = -25;
assign rom[379][1] = -23;
assign rom[379][2] = 9;
assign rom[379][3] = -2;
assign rom[379][4] = 23;
assign rom[379][5] = -26;
assign rom[379][6] = -3;
assign rom[379][7] = 18;
assign rom[379][8] = -9;
assign rom[379][9] = 22;
assign rom[380][0] = -6;
assign rom[380][1] = -32;
assign rom[380][2] = -13;
assign rom[380][3] = -7;
assign rom[380][4] = 29;
assign rom[380][5] = -15;
assign rom[380][6] = -9;
assign rom[380][7] = 22;
assign rom[380][8] = -16;
assign rom[380][9] = 4;
assign rom[381][0] = -8;
assign rom[381][1] = -43;
assign rom[381][2] = -15;
assign rom[381][3] = 3;
assign rom[381][4] = 16;
assign rom[381][5] = -10;
assign rom[381][6] = -9;
assign rom[381][7] = 16;
assign rom[381][8] = -22;
assign rom[381][9] = 6;
assign rom[382][0] = 2;
assign rom[382][1] = -34;
assign rom[382][2] = -14;
assign rom[382][3] = 4;
assign rom[382][4] = 10;
assign rom[382][5] = -8;
assign rom[382][6] = -11;
assign rom[382][7] = 21;
assign rom[382][8] = -20;
assign rom[382][9] = -11;
assign rom[383][0] = -4;
assign rom[383][1] = -27;
assign rom[383][2] = -3;
assign rom[383][3] = 7;
assign rom[383][4] = 3;
assign rom[383][5] = 0;
assign rom[383][6] = -5;
assign rom[383][7] = 20;
assign rom[383][8] = -30;
assign rom[383][9] = -20;
assign rom[384][0] = 16;
assign rom[384][1] = -20;
assign rom[384][2] = -5;
assign rom[384][3] = 2;
assign rom[384][4] = 10;
assign rom[384][5] = -7;
assign rom[384][6] = 5;
assign rom[384][7] = 22;
assign rom[384][8] = -23;
assign rom[384][9] = -16;
assign rom[385][0] = 23;
assign rom[385][1] = -10;
assign rom[385][2] = -18;
assign rom[385][3] = 3;
assign rom[385][4] = -6;
assign rom[385][5] = -1;
assign rom[385][6] = 6;
assign rom[385][7] = 14;
assign rom[385][8] = -25;
assign rom[385][9] = -33;
assign rom[386][0] = 21;
assign rom[386][1] = -10;
assign rom[386][2] = 8;
assign rom[386][3] = 1;
assign rom[386][4] = 1;
assign rom[386][5] = -13;
assign rom[386][6] = 17;
assign rom[386][7] = 12;
assign rom[386][8] = -30;
assign rom[386][9] = -40;
assign rom[387][0] = 11;
assign rom[387][1] = 8;
assign rom[387][2] = 25;
assign rom[387][3] = -14;
assign rom[387][4] = -7;
assign rom[387][5] = -5;
assign rom[387][6] = 2;
assign rom[387][7] = -4;
assign rom[387][8] = -12;
assign rom[387][9] = -35;
assign rom[388][0] = -4;
assign rom[388][1] = 9;
assign rom[388][2] = 35;
assign rom[388][3] = -4;
assign rom[388][4] = -13;
assign rom[388][5] = 9;
assign rom[388][6] = -17;
assign rom[388][7] = 3;
assign rom[388][8] = -26;
assign rom[388][9] = -22;
assign rom[389][0] = -16;
assign rom[389][1] = 19;
assign rom[389][2] = 22;
assign rom[389][3] = -20;
assign rom[389][4] = 3;
assign rom[389][5] = 18;
assign rom[389][6] = -11;
assign rom[389][7] = 12;
assign rom[389][8] = -31;
assign rom[389][9] = -3;
assign rom[390][0] = -16;
assign rom[390][1] = 24;
assign rom[390][2] = -16;
assign rom[390][3] = 5;
assign rom[390][4] = 12;
assign rom[390][5] = 10;
assign rom[390][6] = -9;
assign rom[390][7] = 9;
assign rom[390][8] = -31;
assign rom[390][9] = -7;
assign rom[391][0] = -22;
assign rom[391][1] = 12;
assign rom[391][2] = -2;
assign rom[391][3] = 10;
assign rom[391][4] = 0;
assign rom[391][5] = 11;
assign rom[391][6] = -16;
assign rom[391][7] = 5;
assign rom[391][8] = -18;
assign rom[391][9] = -3;
assign rom[392][0] = -4;
assign rom[392][1] = 2;
assign rom[392][2] = 11;
assign rom[392][3] = 23;
assign rom[392][4] = -6;
assign rom[392][5] = 8;
assign rom[392][6] = -32;
assign rom[392][7] = 0;
assign rom[392][8] = -21;
assign rom[392][9] = -8;
assign rom[393][0] = 10;
assign rom[393][1] = -8;
assign rom[393][2] = 17;
assign rom[393][3] = 16;
assign rom[393][4] = 0;
assign rom[393][5] = -9;
assign rom[393][6] = -16;
assign rom[393][7] = -7;
assign rom[393][8] = -31;
assign rom[393][9] = -7;
assign rom[394][0] = 10;
assign rom[394][1] = -24;
assign rom[394][2] = 5;
assign rom[394][3] = -5;
assign rom[394][4] = 9;
assign rom[394][5] = -4;
assign rom[394][6] = 1;
assign rom[394][7] = -8;
assign rom[394][8] = -36;
assign rom[394][9] = -10;
assign rom[395][0] = 12;
assign rom[395][1] = -39;
assign rom[395][2] = 16;
assign rom[395][3] = -15;
assign rom[395][4] = 30;
assign rom[395][5] = -19;
assign rom[395][6] = 4;
assign rom[395][7] = -12;
assign rom[395][8] = -14;
assign rom[395][9] = -7;
assign rom[396][0] = 8;
assign rom[396][1] = -28;
assign rom[396][2] = 4;
assign rom[396][3] = -19;
assign rom[396][4] = 20;
assign rom[396][5] = -39;
assign rom[396][6] = 10;
assign rom[396][7] = -8;
assign rom[396][8] = -6;
assign rom[396][9] = 0;
assign rom[397][0] = 19;
assign rom[397][1] = -16;
assign rom[397][2] = 11;
assign rom[397][3] = -32;
assign rom[397][4] = 28;
assign rom[397][5] = -30;
assign rom[397][6] = 4;
assign rom[397][7] = -13;
assign rom[397][8] = 1;
assign rom[397][9] = 5;
assign rom[398][0] = 24;
assign rom[398][1] = -16;
assign rom[398][2] = -1;
assign rom[398][3] = -43;
assign rom[398][4] = 8;
assign rom[398][5] = -19;
assign rom[398][6] = 29;
assign rom[398][7] = -30;
assign rom[398][8] = -4;
assign rom[398][9] = 19;
assign rom[399][0] = 11;
assign rom[399][1] = -19;
assign rom[399][2] = 3;
assign rom[399][3] = -38;
assign rom[399][4] = 2;
assign rom[399][5] = -18;
assign rom[399][6] = 26;
assign rom[399][7] = -32;
assign rom[399][8] = 19;
assign rom[399][9] = 17;
assign rom[400][0] = -6;
assign rom[400][1] = 0;
assign rom[400][2] = 11;
assign rom[400][3] = -30;
assign rom[400][4] = -1;
assign rom[400][5] = -27;
assign rom[400][6] = 20;
assign rom[400][7] = -33;
assign rom[400][8] = 17;
assign rom[400][9] = 0;
assign rom[401][0] = -44;
assign rom[401][1] = 19;
assign rom[401][2] = 23;
assign rom[401][3] = -13;
assign rom[401][4] = 6;
assign rom[401][5] = -24;
assign rom[401][6] = 3;
assign rom[401][7] = -29;
assign rom[401][8] = 29;
assign rom[401][9] = -7;
assign rom[402][0] = -63;
assign rom[402][1] = 37;
assign rom[402][2] = 19;
assign rom[402][3] = -11;
assign rom[402][4] = 14;
assign rom[402][5] = -32;
assign rom[402][6] = 7;
assign rom[402][7] = 2;
assign rom[402][8] = 10;
assign rom[402][9] = -17;
assign rom[403][0] = -62;
assign rom[403][1] = 24;
assign rom[403][2] = 13;
assign rom[403][3] = -10;
assign rom[403][4] = 28;
assign rom[403][5] = -14;
assign rom[403][6] = 4;
assign rom[403][7] = -2;
assign rom[403][8] = 0;
assign rom[403][9] = -5;
assign rom[404][0] = -36;
assign rom[404][1] = -3;
assign rom[404][2] = 14;
assign rom[404][3] = -8;
assign rom[404][4] = 28;
assign rom[404][5] = -12;
assign rom[404][6] = -5;
assign rom[404][7] = 3;
assign rom[404][8] = 7;
assign rom[404][9] = 12;
assign rom[405][0] = -24;
assign rom[405][1] = -27;
assign rom[405][2] = 6;
assign rom[405][3] = 3;
assign rom[405][4] = 37;
assign rom[405][5] = -12;
assign rom[405][6] = -8;
assign rom[405][7] = 14;
assign rom[405][8] = 4;
assign rom[405][9] = 21;
assign rom[406][0] = -4;
assign rom[406][1] = -38;
assign rom[406][2] = -8;
assign rom[406][3] = -4;
assign rom[406][4] = 19;
assign rom[406][5] = -7;
assign rom[406][6] = -5;
assign rom[406][7] = 5;
assign rom[406][8] = -13;
assign rom[406][9] = 5;
assign rom[407][0] = -4;
assign rom[407][1] = -40;
assign rom[407][2] = -10;
assign rom[407][3] = 1;
assign rom[407][4] = 12;
assign rom[407][5] = -8;
assign rom[407][6] = -6;
assign rom[407][7] = 10;
assign rom[407][8] = -24;
assign rom[407][9] = -12;
assign rom[408][0] = 4;
assign rom[408][1] = -43;
assign rom[408][2] = 1;
assign rom[408][3] = 10;
assign rom[408][4] = 13;
assign rom[408][5] = -6;
assign rom[408][6] = 5;
assign rom[408][7] = 23;
assign rom[408][8] = -21;
assign rom[408][9] = -6;
assign rom[409][0] = -2;
assign rom[409][1] = -26;
assign rom[409][2] = 7;
assign rom[409][3] = 13;
assign rom[409][4] = -7;
assign rom[409][5] = 6;
assign rom[409][6] = -4;
assign rom[409][7] = 13;
assign rom[409][8] = -18;
assign rom[409][9] = -20;
assign rom[410][0] = 2;
assign rom[410][1] = -26;
assign rom[410][2] = -2;
assign rom[410][3] = 23;
assign rom[410][4] = 2;
assign rom[410][5] = 5;
assign rom[410][6] = -6;
assign rom[410][7] = 4;
assign rom[410][8] = -27;
assign rom[410][9] = -30;
assign rom[411][0] = 21;
assign rom[411][1] = -24;
assign rom[411][2] = 3;
assign rom[411][3] = 11;
assign rom[411][4] = -17;
assign rom[411][5] = -4;
assign rom[411][6] = -6;
assign rom[411][7] = 7;
assign rom[411][8] = -11;
assign rom[411][9] = -32;
assign rom[412][0] = 15;
assign rom[412][1] = -17;
assign rom[412][2] = 14;
assign rom[412][3] = 5;
assign rom[412][4] = -13;
assign rom[412][5] = -6;
assign rom[412][6] = 1;
assign rom[412][7] = 3;
assign rom[412][8] = -20;
assign rom[412][9] = -40;
assign rom[413][0] = 1;
assign rom[413][1] = 1;
assign rom[413][2] = 31;
assign rom[413][3] = -14;
assign rom[413][4] = -18;
assign rom[413][5] = 9;
assign rom[413][6] = -3;
assign rom[413][7] = -13;
assign rom[413][8] = -22;
assign rom[413][9] = -36;
assign rom[414][0] = -3;
assign rom[414][1] = 12;
assign rom[414][2] = 47;
assign rom[414][3] = -8;
assign rom[414][4] = -21;
assign rom[414][5] = 6;
assign rom[414][6] = -19;
assign rom[414][7] = 10;
assign rom[414][8] = -21;
assign rom[414][9] = -19;
assign rom[415][0] = -18;
assign rom[415][1] = 20;
assign rom[415][2] = 33;
assign rom[415][3] = -14;
assign rom[415][4] = 8;
assign rom[415][5] = 11;
assign rom[415][6] = -13;
assign rom[415][7] = 12;
assign rom[415][8] = -32;
assign rom[415][9] = -14;
assign rom[416][0] = -6;
assign rom[416][1] = 22;
assign rom[416][2] = -2;
assign rom[416][3] = 1;
assign rom[416][4] = -1;
assign rom[416][5] = 15;
assign rom[416][6] = 0;
assign rom[416][7] = 9;
assign rom[416][8] = -17;
assign rom[416][9] = 4;
assign rom[417][0] = -19;
assign rom[417][1] = 15;
assign rom[417][2] = 7;
assign rom[417][3] = 27;
assign rom[417][4] = -10;
assign rom[417][5] = 7;
assign rom[417][6] = -15;
assign rom[417][7] = 5;
assign rom[417][8] = -25;
assign rom[417][9] = -7;
assign rom[418][0] = -17;
assign rom[418][1] = 15;
assign rom[418][2] = 6;
assign rom[418][3] = 25;
assign rom[418][4] = -23;
assign rom[418][5] = 9;
assign rom[418][6] = -26;
assign rom[418][7] = -2;
assign rom[418][8] = -22;
assign rom[418][9] = -14;
assign rom[419][0] = 1;
assign rom[419][1] = -18;
assign rom[419][2] = 20;
assign rom[419][3] = 27;
assign rom[419][4] = -12;
assign rom[419][5] = 1;
assign rom[419][6] = -31;
assign rom[419][7] = -11;
assign rom[419][8] = -30;
assign rom[419][9] = -9;
assign rom[420][0] = 15;
assign rom[420][1] = -36;
assign rom[420][2] = 17;
assign rom[420][3] = 1;
assign rom[420][4] = -6;
assign rom[420][5] = 20;
assign rom[420][6] = -14;
assign rom[420][7] = -15;
assign rom[420][8] = -19;
assign rom[420][9] = -11;
assign rom[421][0] = 7;
assign rom[421][1] = -35;
assign rom[421][2] = 22;
assign rom[421][3] = -9;
assign rom[421][4] = -3;
assign rom[421][5] = 9;
assign rom[421][6] = -8;
assign rom[421][7] = -22;
assign rom[421][8] = -6;
assign rom[421][9] = -1;
assign rom[422][0] = 9;
assign rom[422][1] = -21;
assign rom[422][2] = 3;
assign rom[422][3] = -16;
assign rom[422][4] = 19;
assign rom[422][5] = -21;
assign rom[422][6] = 10;
assign rom[422][7] = -14;
assign rom[422][8] = 11;
assign rom[422][9] = 9;
assign rom[423][0] = 7;
assign rom[423][1] = -16;
assign rom[423][2] = 12;
assign rom[423][3] = -36;
assign rom[423][4] = 17;
assign rom[423][5] = -34;
assign rom[423][6] = 1;
assign rom[423][7] = -22;
assign rom[423][8] = 12;
assign rom[423][9] = 5;
assign rom[424][0] = 17;
assign rom[424][1] = -16;
assign rom[424][2] = 1;
assign rom[424][3] = -50;
assign rom[424][4] = 0;
assign rom[424][5] = -32;
assign rom[424][6] = 22;
assign rom[424][7] = -26;
assign rom[424][8] = 24;
assign rom[424][9] = 5;
assign rom[425][0] = 10;
assign rom[425][1] = 3;
assign rom[425][2] = 16;
assign rom[425][3] = -40;
assign rom[425][4] = -9;
assign rom[425][5] = -41;
assign rom[425][6] = 32;
assign rom[425][7] = -27;
assign rom[425][8] = 19;
assign rom[425][9] = 13;
assign rom[426][0] = -11;
assign rom[426][1] = 10;
assign rom[426][2] = 26;
assign rom[426][3] = -35;
assign rom[426][4] = 5;
assign rom[426][5] = -31;
assign rom[426][6] = 22;
assign rom[426][7] = -17;
assign rom[426][8] = 27;
assign rom[426][9] = 5;
assign rom[427][0] = -48;
assign rom[427][1] = 18;
assign rom[427][2] = 20;
assign rom[427][3] = -38;
assign rom[427][4] = 9;
assign rom[427][5] = -24;
assign rom[427][6] = 15;
assign rom[427][7] = 2;
assign rom[427][8] = 18;
assign rom[427][9] = -11;
assign rom[428][0] = -59;
assign rom[428][1] = 36;
assign rom[428][2] = 16;
assign rom[428][3] = -37;
assign rom[428][4] = 25;
assign rom[428][5] = -24;
assign rom[428][6] = 4;
assign rom[428][7] = 0;
assign rom[428][8] = 3;
assign rom[428][9] = -18;
assign rom[429][0] = -44;
assign rom[429][1] = 25;
assign rom[429][2] = 8;
assign rom[429][3] = -22;
assign rom[429][4] = 30;
assign rom[429][5] = -22;
assign rom[429][6] = -4;
assign rom[429][7] = 14;
assign rom[429][8] = -10;
assign rom[429][9] = 1;
assign rom[430][0] = -20;
assign rom[430][1] = -11;
assign rom[430][2] = 5;
assign rom[430][3] = -3;
assign rom[430][4] = 33;
assign rom[430][5] = 0;
assign rom[430][6] = -10;
assign rom[430][7] = 5;
assign rom[430][8] = 1;
assign rom[430][9] = 5;
assign rom[431][0] = -10;
assign rom[431][1] = -26;
assign rom[431][2] = 3;
assign rom[431][3] = 4;
assign rom[431][4] = 29;
assign rom[431][5] = 0;
assign rom[431][6] = 4;
assign rom[431][7] = -9;
assign rom[431][8] = -2;
assign rom[431][9] = 1;
assign rom[432][0] = 6;
assign rom[432][1] = -39;
assign rom[432][2] = 8;
assign rom[432][3] = 17;
assign rom[432][4] = 8;
assign rom[432][5] = 8;
assign rom[432][6] = -6;
assign rom[432][7] = 4;
assign rom[432][8] = -4;
assign rom[432][9] = -9;
assign rom[433][0] = 7;
assign rom[433][1] = -42;
assign rom[433][2] = 0;
assign rom[433][3] = 17;
assign rom[433][4] = -6;
assign rom[433][5] = -6;
assign rom[433][6] = 11;
assign rom[433][7] = 13;
assign rom[433][8] = -22;
assign rom[433][9] = -5;
assign rom[434][0] = -4;
assign rom[434][1] = -24;
assign rom[434][2] = 8;
assign rom[434][3] = 19;
assign rom[434][4] = -5;
assign rom[434][5] = 10;
assign rom[434][6] = 5;
assign rom[434][7] = 3;
assign rom[434][8] = -14;
assign rom[434][9] = -13;
assign rom[435][0] = 6;
assign rom[435][1] = -10;
assign rom[435][2] = 11;
assign rom[435][3] = 24;
assign rom[435][4] = -6;
assign rom[435][5] = 9;
assign rom[435][6] = 8;
assign rom[435][7] = 4;
assign rom[435][8] = -9;
assign rom[435][9] = -18;
assign rom[436][0] = 2;
assign rom[436][1] = -17;
assign rom[436][2] = 10;
assign rom[436][3] = 22;
assign rom[436][4] = -16;
assign rom[436][5] = 1;
assign rom[436][6] = 0;
assign rom[436][7] = -8;
assign rom[436][8] = -23;
assign rom[436][9] = -31;
assign rom[437][0] = 12;
assign rom[437][1] = -11;
assign rom[437][2] = 24;
assign rom[437][3] = 17;
assign rom[437][4] = -31;
assign rom[437][5] = 6;
assign rom[437][6] = 1;
assign rom[437][7] = -21;
assign rom[437][8] = -1;
assign rom[437][9] = -38;
assign rom[438][0] = -2;
assign rom[438][1] = -18;
assign rom[438][2] = 23;
assign rom[438][3] = 5;
assign rom[438][4] = -22;
assign rom[438][5] = 11;
assign rom[438][6] = -8;
assign rom[438][7] = -9;
assign rom[438][8] = -4;
assign rom[438][9] = -38;
assign rom[439][0] = 1;
assign rom[439][1] = 0;
assign rom[439][2] = 49;
assign rom[439][3] = -11;
assign rom[439][4] = -26;
assign rom[439][5] = 3;
assign rom[439][6] = -27;
assign rom[439][7] = -11;
assign rom[439][8] = -9;
assign rom[439][9] = -25;
assign rom[440][0] = -4;
assign rom[440][1] = 15;
assign rom[440][2] = 45;
assign rom[440][3] = -23;
assign rom[440][4] = -16;
assign rom[440][5] = 19;
assign rom[440][6] = -19;
assign rom[440][7] = 3;
assign rom[440][8] = -31;
assign rom[440][9] = -8;
assign rom[441][0] = -9;
assign rom[441][1] = 21;
assign rom[441][2] = 23;
assign rom[441][3] = -6;
assign rom[441][4] = 7;
assign rom[441][5] = 4;
assign rom[441][6] = -15;
assign rom[441][7] = 12;
assign rom[441][8] = -28;
assign rom[441][9] = -12;
assign rom[442][0] = -1;
assign rom[442][1] = 24;
assign rom[442][2] = -2;
assign rom[442][3] = 11;
assign rom[442][4] = 8;
assign rom[442][5] = 16;
assign rom[442][6] = -11;
assign rom[442][7] = 19;
assign rom[442][8] = -20;
assign rom[442][9] = -10;
assign rom[443][0] = -23;
assign rom[443][1] = 20;
assign rom[443][2] = -9;
assign rom[443][3] = 21;
assign rom[443][4] = 3;
assign rom[443][5] = 12;
assign rom[443][6] = -16;
assign rom[443][7] = -6;
assign rom[443][8] = -27;
assign rom[443][9] = -18;
assign rom[444][0] = -16;
assign rom[444][1] = 4;
assign rom[444][2] = 17;
assign rom[444][3] = 38;
assign rom[444][4] = -18;
assign rom[444][5] = 13;
assign rom[444][6] = -39;
assign rom[444][7] = -10;
assign rom[444][8] = -23;
assign rom[444][9] = -17;
assign rom[445][0] = -5;
assign rom[445][1] = -27;
assign rom[445][2] = 21;
assign rom[445][3] = 32;
assign rom[445][4] = -24;
assign rom[445][5] = 3;
assign rom[445][6] = -30;
assign rom[445][7] = -11;
assign rom[445][8] = -21;
assign rom[445][9] = -23;
assign rom[446][0] = 2;
assign rom[446][1] = -37;
assign rom[446][2] = 21;
assign rom[446][3] = 29;
assign rom[446][4] = -22;
assign rom[446][5] = 28;
assign rom[446][6] = -23;
assign rom[446][7] = -17;
assign rom[446][8] = -14;
assign rom[446][9] = -14;
assign rom[447][0] = 16;
assign rom[447][1] = -32;
assign rom[447][2] = 21;
assign rom[447][3] = 17;
assign rom[447][4] = -18;
assign rom[447][5] = 32;
assign rom[447][6] = -18;
assign rom[447][7] = -39;
assign rom[447][8] = 3;
assign rom[447][9] = -19;
assign rom[448][0] = 19;
assign rom[448][1] = -29;
assign rom[448][2] = 14;
assign rom[448][3] = 0;
assign rom[448][4] = -20;
assign rom[448][5] = 9;
assign rom[448][6] = -6;
assign rom[448][7] = -36;
assign rom[448][8] = 4;
assign rom[448][9] = -5;
assign rom[449][0] = 18;
assign rom[449][1] = -15;
assign rom[449][2] = 11;
assign rom[449][3] = -19;
assign rom[449][4] = -12;
assign rom[449][5] = -14;
assign rom[449][6] = 2;
assign rom[449][7] = -27;
assign rom[449][8] = 18;
assign rom[449][9] = -9;
assign rom[450][0] = 13;
assign rom[450][1] = -9;
assign rom[450][2] = 7;
assign rom[450][3] = -39;
assign rom[450][4] = -20;
assign rom[450][5] = -30;
assign rom[450][6] = 11;
assign rom[450][7] = -46;
assign rom[450][8] = 19;
assign rom[450][9] = 0;
assign rom[451][0] = 9;
assign rom[451][1] = -1;
assign rom[451][2] = 14;
assign rom[451][3] = -38;
assign rom[451][4] = -17;
assign rom[451][5] = -34;
assign rom[451][6] = 30;
assign rom[451][7] = -22;
assign rom[451][8] = 17;
assign rom[451][9] = 0;
assign rom[452][0] = -5;
assign rom[452][1] = 9;
assign rom[452][2] = 24;
assign rom[452][3] = -39;
assign rom[452][4] = -7;
assign rom[452][5] = -18;
assign rom[452][6] = 31;
assign rom[452][7] = -20;
assign rom[452][8] = 8;
assign rom[452][9] = -8;
assign rom[453][0] = -18;
assign rom[453][1] = 11;
assign rom[453][2] = 15;
assign rom[453][3] = -44;
assign rom[453][4] = -1;
assign rom[453][5] = -16;
assign rom[453][6] = 7;
assign rom[453][7] = 10;
assign rom[453][8] = 4;
assign rom[453][9] = -11;
assign rom[454][0] = -30;
assign rom[454][1] = 17;
assign rom[454][2] = 23;
assign rom[454][3] = -38;
assign rom[454][4] = 11;
assign rom[454][5] = -6;
assign rom[454][6] = 9;
assign rom[454][7] = 14;
assign rom[454][8] = -8;
assign rom[454][9] = -9;
assign rom[455][0] = -27;
assign rom[455][1] = 18;
assign rom[455][2] = 13;
assign rom[455][3] = -27;
assign rom[455][4] = 14;
assign rom[455][5] = 7;
assign rom[455][6] = 12;
assign rom[455][7] = 3;
assign rom[455][8] = -5;
assign rom[455][9] = 2;
assign rom[456][0] = -15;
assign rom[456][1] = -4;
assign rom[456][2] = 14;
assign rom[456][3] = -4;
assign rom[456][4] = 14;
assign rom[456][5] = -9;
assign rom[456][6] = 3;
assign rom[456][7] = -10;
assign rom[456][8] = -5;
assign rom[456][9] = 4;
assign rom[457][0] = 4;
assign rom[457][1] = -22;
assign rom[457][2] = 17;
assign rom[457][3] = 9;
assign rom[457][4] = -2;
assign rom[457][5] = 6;
assign rom[457][6] = 13;
assign rom[457][7] = -5;
assign rom[457][8] = -7;
assign rom[457][9] = -7;
assign rom[458][0] = 6;
assign rom[458][1] = -32;
assign rom[458][2] = 9;
assign rom[458][3] = 19;
assign rom[458][4] = -12;
assign rom[458][5] = 13;
assign rom[458][6] = 19;
assign rom[458][7] = -18;
assign rom[458][8] = -13;
assign rom[458][9] = -9;
assign rom[459][0] = 8;
assign rom[459][1] = -17;
assign rom[459][2] = 11;
assign rom[459][3] = 13;
assign rom[459][4] = -15;
assign rom[459][5] = 9;
assign rom[459][6] = 12;
assign rom[459][7] = -14;
assign rom[459][8] = -10;
assign rom[459][9] = -20;
assign rom[460][0] = -3;
assign rom[460][1] = -9;
assign rom[460][2] = 6;
assign rom[460][3] = 19;
assign rom[460][4] = -27;
assign rom[460][5] = 1;
assign rom[460][6] = 15;
assign rom[460][7] = -26;
assign rom[460][8] = -2;
assign rom[460][9] = -14;
assign rom[461][0] = 1;
assign rom[461][1] = -10;
assign rom[461][2] = 2;
assign rom[461][3] = 11;
assign rom[461][4] = -18;
assign rom[461][5] = 3;
assign rom[461][6] = -5;
assign rom[461][7] = -18;
assign rom[461][8] = -7;
assign rom[461][9] = -18;
assign rom[462][0] = 9;
assign rom[462][1] = -23;
assign rom[462][2] = 10;
assign rom[462][3] = 8;
assign rom[462][4] = -23;
assign rom[462][5] = 1;
assign rom[462][6] = 6;
assign rom[462][7] = -29;
assign rom[462][8] = -3;
assign rom[462][9] = -16;
assign rom[463][0] = 6;
assign rom[463][1] = -29;
assign rom[463][2] = 19;
assign rom[463][3] = 12;
assign rom[463][4] = -26;
assign rom[463][5] = 6;
assign rom[463][6] = 0;
assign rom[463][7] = -39;
assign rom[463][8] = -4;
assign rom[463][9] = -32;
assign rom[464][0] = 0;
assign rom[464][1] = -6;
assign rom[464][2] = 32;
assign rom[464][3] = -3;
assign rom[464][4] = -32;
assign rom[464][5] = 2;
assign rom[464][6] = -22;
assign rom[464][7] = -22;
assign rom[464][8] = -15;
assign rom[464][9] = -33;
assign rom[465][0] = -16;
assign rom[465][1] = -11;
assign rom[465][2] = 36;
assign rom[465][3] = -17;
assign rom[465][4] = -21;
assign rom[465][5] = 9;
assign rom[465][6] = -11;
assign rom[465][7] = -17;
assign rom[465][8] = -11;
assign rom[465][9] = -33;
assign rom[466][0] = -8;
assign rom[466][1] = 12;
assign rom[466][2] = 36;
assign rom[466][3] = -15;
assign rom[466][4] = 0;
assign rom[466][5] = 19;
assign rom[466][6] = -23;
assign rom[466][7] = 8;
assign rom[466][8] = -19;
assign rom[466][9] = -5;
assign rom[467][0] = -13;
assign rom[467][1] = 16;
assign rom[467][2] = 20;
assign rom[467][3] = -23;
assign rom[467][4] = -2;
assign rom[467][5] = 20;
assign rom[467][6] = -10;
assign rom[467][7] = 12;
assign rom[467][8] = -30;
assign rom[467][9] = -8;
assign rom[468][0] = -10;
assign rom[468][1] = 11;
assign rom[468][2] = -10;
assign rom[468][3] = -6;
assign rom[468][4] = 1;
assign rom[468][5] = 13;
assign rom[468][6] = 0;
assign rom[468][7] = 5;
assign rom[468][8] = -33;
assign rom[468][9] = -10;
assign rom[469][0] = -30;
assign rom[469][1] = 15;
assign rom[469][2] = -2;
assign rom[469][3] = 21;
assign rom[469][4] = -12;
assign rom[469][5] = 0;
assign rom[469][6] = -10;
assign rom[469][7] = 2;
assign rom[469][8] = -37;
assign rom[469][9] = -16;
assign rom[470][0] = -17;
assign rom[470][1] = -4;
assign rom[470][2] = 0;
assign rom[470][3] = 29;
assign rom[470][4] = -9;
assign rom[470][5] = 2;
assign rom[470][6] = -36;
assign rom[470][7] = -18;
assign rom[470][8] = -25;
assign rom[470][9] = -12;
assign rom[471][0] = 3;
assign rom[471][1] = -23;
assign rom[471][2] = 11;
assign rom[471][3] = 42;
assign rom[471][4] = -22;
assign rom[471][5] = 12;
assign rom[471][6] = -26;
assign rom[471][7] = -13;
assign rom[471][8] = -19;
assign rom[471][9] = -24;
assign rom[472][0] = 13;
assign rom[472][1] = -32;
assign rom[472][2] = 22;
assign rom[472][3] = 29;
assign rom[472][4] = -21;
assign rom[472][5] = 24;
assign rom[472][6] = -23;
assign rom[472][7] = -27;
assign rom[472][8] = -14;
assign rom[472][9] = -22;
assign rom[473][0] = 4;
assign rom[473][1] = -22;
assign rom[473][2] = 23;
assign rom[473][3] = 11;
assign rom[473][4] = -28;
assign rom[473][5] = 20;
assign rom[473][6] = -14;
assign rom[473][7] = -35;
assign rom[473][8] = 3;
assign rom[473][9] = -32;
assign rom[474][0] = 3;
assign rom[474][1] = -20;
assign rom[474][2] = 12;
assign rom[474][3] = 13;
assign rom[474][4] = -41;
assign rom[474][5] = 21;
assign rom[474][6] = -8;
assign rom[474][7] = -30;
assign rom[474][8] = 2;
assign rom[474][9] = -19;
assign rom[475][0] = 16;
assign rom[475][1] = -9;
assign rom[475][2] = 20;
assign rom[475][3] = 6;
assign rom[475][4] = -31;
assign rom[475][5] = 14;
assign rom[475][6] = 11;
assign rom[475][7] = -30;
assign rom[475][8] = 9;
assign rom[475][9] = -16;
assign rom[476][0] = 13;
assign rom[476][1] = -2;
assign rom[476][2] = 21;
assign rom[476][3] = -8;
assign rom[476][4] = -47;
assign rom[476][5] = 4;
assign rom[476][6] = 18;
assign rom[476][7] = -24;
assign rom[476][8] = 3;
assign rom[476][9] = -27;
assign rom[477][0] = 15;
assign rom[477][1] = 1;
assign rom[477][2] = 17;
assign rom[477][3] = -15;
assign rom[477][4] = -32;
assign rom[477][5] = 7;
assign rom[477][6] = 28;
assign rom[477][7] = -16;
assign rom[477][8] = -4;
assign rom[477][9] = -25;
assign rom[478][0] = 17;
assign rom[478][1] = -1;
assign rom[478][2] = 8;
assign rom[478][3] = -29;
assign rom[478][4] = -33;
assign rom[478][5] = 0;
assign rom[478][6] = 28;
assign rom[478][7] = -10;
assign rom[478][8] = -8;
assign rom[478][9] = -33;
assign rom[479][0] = 3;
assign rom[479][1] = 10;
assign rom[479][2] = 14;
assign rom[479][3] = -19;
assign rom[479][4] = -16;
assign rom[479][5] = -4;
assign rom[479][6] = 27;
assign rom[479][7] = 0;
assign rom[479][8] = -7;
assign rom[479][9] = -18;
assign rom[480][0] = -17;
assign rom[480][1] = 11;
assign rom[480][2] = 5;
assign rom[480][3] = -15;
assign rom[480][4] = -6;
assign rom[480][5] = -2;
assign rom[480][6] = 26;
assign rom[480][7] = -1;
assign rom[480][8] = -18;
assign rom[480][9] = -4;
assign rom[481][0] = -13;
assign rom[481][1] = 1;
assign rom[481][2] = 13;
assign rom[481][3] = -9;
assign rom[481][4] = 1;
assign rom[481][5] = 3;
assign rom[481][6] = 14;
assign rom[481][7] = 5;
assign rom[481][8] = -9;
assign rom[481][9] = -9;
assign rom[482][0] = 0;
assign rom[482][1] = -21;
assign rom[482][2] = 4;
assign rom[482][3] = -3;
assign rom[482][4] = -3;
assign rom[482][5] = -3;
assign rom[482][6] = 21;
assign rom[482][7] = -8;
assign rom[482][8] = -18;
assign rom[482][9] = -4;
assign rom[483][0] = -1;
assign rom[483][1] = -17;
assign rom[483][2] = 8;
assign rom[483][3] = 10;
assign rom[483][4] = -4;
assign rom[483][5] = -5;
assign rom[483][6] = 29;
assign rom[483][7] = -22;
assign rom[483][8] = -15;
assign rom[483][9] = -6;
assign rom[484][0] = 2;
assign rom[484][1] = -4;
assign rom[484][2] = 15;
assign rom[484][3] = 23;
assign rom[484][4] = -13;
assign rom[484][5] = 9;
assign rom[484][6] = 14;
assign rom[484][7] = -21;
assign rom[484][8] = -4;
assign rom[484][9] = -15;
assign rom[485][0] = -6;
assign rom[485][1] = 0;
assign rom[485][2] = 14;
assign rom[485][3] = 28;
assign rom[485][4] = -8;
assign rom[485][5] = 1;
assign rom[485][6] = 17;
assign rom[485][7] = -19;
assign rom[485][8] = 1;
assign rom[485][9] = -22;
assign rom[486][0] = -9;
assign rom[486][1] = -6;
assign rom[486][2] = 13;
assign rom[486][3] = 16;
assign rom[486][4] = -16;
assign rom[486][5] = 3;
assign rom[486][6] = 16;
assign rom[486][7] = -27;
assign rom[486][8] = 2;
assign rom[486][9] = -5;
assign rom[487][0] = -10;
assign rom[487][1] = -19;
assign rom[487][2] = 3;
assign rom[487][3] = 5;
assign rom[487][4] = -25;
assign rom[487][5] = 14;
assign rom[487][6] = 6;
assign rom[487][7] = -49;
assign rom[487][8] = -8;
assign rom[487][9] = -1;
assign rom[488][0] = 5;
assign rom[488][1] = -27;
assign rom[488][2] = 15;
assign rom[488][3] = 15;
assign rom[488][4] = -26;
assign rom[488][5] = -3;
assign rom[488][6] = -12;
assign rom[488][7] = -44;
assign rom[488][8] = 2;
assign rom[488][9] = -20;
assign rom[489][0] = -7;
assign rom[489][1] = -11;
assign rom[489][2] = 19;
assign rom[489][3] = -3;
assign rom[489][4] = -23;
assign rom[489][5] = 16;
assign rom[489][6] = -1;
assign rom[489][7] = -31;
assign rom[489][8] = 7;
assign rom[489][9] = -11;
assign rom[490][0] = -11;
assign rom[490][1] = -13;
assign rom[490][2] = 39;
assign rom[490][3] = -21;
assign rom[490][4] = -20;
assign rom[490][5] = 16;
assign rom[490][6] = -13;
assign rom[490][7] = -28;
assign rom[490][8] = -13;
assign rom[490][9] = -22;
assign rom[491][0] = -21;
assign rom[491][1] = 0;
assign rom[491][2] = 30;
assign rom[491][3] = -31;
assign rom[491][4] = -10;
assign rom[491][5] = 19;
assign rom[491][6] = -24;
assign rom[491][7] = -7;
assign rom[491][8] = -18;
assign rom[491][9] = -13;
assign rom[492][0] = -10;
assign rom[492][1] = 10;
assign rom[492][2] = 28;
assign rom[492][3] = -21;
assign rom[492][4] = -5;
assign rom[492][5] = 19;
assign rom[492][6] = -20;
assign rom[492][7] = -1;
assign rom[492][8] = -32;
assign rom[492][9] = 0;
assign rom[493][0] = -3;
assign rom[493][1] = 28;
assign rom[493][2] = 11;
assign rom[493][3] = -15;
assign rom[493][4] = 8;
assign rom[493][5] = 10;
assign rom[493][6] = -9;
assign rom[493][7] = 11;
assign rom[493][8] = -34;
assign rom[493][9] = -5;
assign rom[494][0] = -15;
assign rom[494][1] = 13;
assign rom[494][2] = 1;
assign rom[494][3] = 3;
assign rom[494][4] = 12;
assign rom[494][5] = 13;
assign rom[494][6] = -3;
assign rom[494][7] = 13;
assign rom[494][8] = -31;
assign rom[494][9] = -3;
assign rom[495][0] = -22;
assign rom[495][1] = 18;
assign rom[495][2] = -5;
assign rom[495][3] = 12;
assign rom[495][4] = -7;
assign rom[495][5] = -8;
assign rom[495][6] = -14;
assign rom[495][7] = -2;
assign rom[495][8] = -25;
assign rom[495][9] = -20;
assign rom[496][0] = -27;
assign rom[496][1] = -1;
assign rom[496][2] = 7;
assign rom[496][3] = 34;
assign rom[496][4] = -24;
assign rom[496][5] = 7;
assign rom[496][6] = -16;
assign rom[496][7] = -21;
assign rom[496][8] = -37;
assign rom[496][9] = -7;
assign rom[497][0] = -4;
assign rom[497][1] = 4;
assign rom[497][2] = 18;
assign rom[497][3] = 24;
assign rom[497][4] = -17;
assign rom[497][5] = -5;
assign rom[497][6] = -39;
assign rom[497][7] = -15;
assign rom[497][8] = -11;
assign rom[497][9] = -15;
assign rom[498][0] = 3;
assign rom[498][1] = -13;
assign rom[498][2] = 17;
assign rom[498][3] = 33;
assign rom[498][4] = -36;
assign rom[498][5] = 3;
assign rom[498][6] = -26;
assign rom[498][7] = -28;
assign rom[498][8] = 7;
assign rom[498][9] = -20;
assign rom[499][0] = -3;
assign rom[499][1] = -7;
assign rom[499][2] = 20;
assign rom[499][3] = 20;
assign rom[499][4] = -39;
assign rom[499][5] = 7;
assign rom[499][6] = -23;
assign rom[499][7] = -23;
assign rom[499][8] = 11;
assign rom[499][9] = -35;
assign rom[500][0] = -4;
assign rom[500][1] = 1;
assign rom[500][2] = 20;
assign rom[500][3] = 11;
assign rom[500][4] = -46;
assign rom[500][5] = 16;
assign rom[500][6] = -23;
assign rom[500][7] = -28;
assign rom[500][8] = 2;
assign rom[500][9] = -32;
assign rom[501][0] = 7;
assign rom[501][1] = 1;
assign rom[501][2] = 17;
assign rom[501][3] = 4;
assign rom[501][4] = -52;
assign rom[501][5] = 16;
assign rom[501][6] = -7;
assign rom[501][7] = -35;
assign rom[501][8] = -2;
assign rom[501][9] = -22;
assign rom[502][0] = 19;
assign rom[502][1] = 7;
assign rom[502][2] = 14;
assign rom[502][3] = 5;
assign rom[502][4] = -37;
assign rom[502][5] = 19;
assign rom[502][6] = 11;
assign rom[502][7] = -13;
assign rom[502][8] = -9;
assign rom[502][9] = -22;
assign rom[503][0] = 18;
assign rom[503][1] = 0;
assign rom[503][2] = 20;
assign rom[503][3] = -12;
assign rom[503][4] = -25;
assign rom[503][5] = 5;
assign rom[503][6] = 18;
assign rom[503][7] = -4;
assign rom[503][8] = -5;
assign rom[503][9] = -40;
assign rom[504][0] = 10;
assign rom[504][1] = -8;
assign rom[504][2] = 17;
assign rom[504][3] = -10;
assign rom[504][4] = -20;
assign rom[504][5] = 4;
assign rom[504][6] = 25;
assign rom[504][7] = -3;
assign rom[504][8] = -21;
assign rom[504][9] = -37;
assign rom[505][0] = 12;
assign rom[505][1] = -1;
assign rom[505][2] = -4;
assign rom[505][3] = -19;
assign rom[505][4] = -11;
assign rom[505][5] = 1;
assign rom[505][6] = 32;
assign rom[505][7] = -1;
assign rom[505][8] = -22;
assign rom[505][9] = -22;
assign rom[506][0] = -5;
assign rom[506][1] = -1;
assign rom[506][2] = -9;
assign rom[506][3] = -7;
assign rom[506][4] = -15;
assign rom[506][5] = -6;
assign rom[506][6] = 30;
assign rom[506][7] = 5;
assign rom[506][8] = -20;
assign rom[506][9] = -6;
assign rom[507][0] = -4;
assign rom[507][1] = -4;
assign rom[507][2] = -9;
assign rom[507][3] = 3;
assign rom[507][4] = -3;
assign rom[507][5] = 5;
assign rom[507][6] = 30;
assign rom[507][7] = -13;
assign rom[507][8] = -2;
assign rom[507][9] = -2;
assign rom[508][0] = 3;
assign rom[508][1] = -12;
assign rom[508][2] = 5;
assign rom[508][3] = 8;
assign rom[508][4] = -1;
assign rom[508][5] = -4;
assign rom[508][6] = 33;
assign rom[508][7] = -21;
assign rom[508][8] = -6;
assign rom[508][9] = -10;
assign rom[509][0] = -2;
assign rom[509][1] = -8;
assign rom[509][2] = -3;
assign rom[509][3] = 10;
assign rom[509][4] = -7;
assign rom[509][5] = 3;
assign rom[509][6] = 22;
assign rom[509][7] = -12;
assign rom[509][8] = -6;
assign rom[509][9] = -12;
assign rom[510][0] = -1;
assign rom[510][1] = -3;
assign rom[510][2] = 9;
assign rom[510][3] = 26;
assign rom[510][4] = -4;
assign rom[510][5] = 12;
assign rom[510][6] = 18;
assign rom[510][7] = -30;
assign rom[510][8] = 0;
assign rom[510][9] = -11;
assign rom[511][0] = -8;
assign rom[511][1] = -3;
assign rom[511][2] = 13;
assign rom[511][3] = 12;
assign rom[511][4] = -17;
assign rom[511][5] = 7;
assign rom[511][6] = 13;
assign rom[511][7] = -35;
assign rom[511][8] = -2;
assign rom[511][9] = -18;
assign rom[512][0] = -3;
assign rom[512][1] = -10;
assign rom[512][2] = 3;
assign rom[512][3] = 4;
assign rom[512][4] = -6;
assign rom[512][5] = 2;
assign rom[512][6] = 8;
assign rom[512][7] = -30;
assign rom[512][8] = -4;
assign rom[512][9] = -21;
assign rom[513][0] = -11;
assign rom[513][1] = -27;
assign rom[513][2] = 5;
assign rom[513][3] = 6;
assign rom[513][4] = -20;
assign rom[513][5] = 0;
assign rom[513][6] = 4;
assign rom[513][7] = -50;
assign rom[513][8] = 2;
assign rom[513][9] = -10;
assign rom[514][0] = -9;
assign rom[514][1] = -14;
assign rom[514][2] = 17;
assign rom[514][3] = -2;
assign rom[514][4] = -25;
assign rom[514][5] = 2;
assign rom[514][6] = -2;
assign rom[514][7] = -48;
assign rom[514][8] = -3;
assign rom[514][9] = -16;
assign rom[515][0] = 1;
assign rom[515][1] = -13;
assign rom[515][2] = 26;
assign rom[515][3] = -10;
assign rom[515][4] = -28;
assign rom[515][5] = 16;
assign rom[515][6] = -19;
assign rom[515][7] = -35;
assign rom[515][8] = 2;
assign rom[515][9] = -20;
assign rom[516][0] = -2;
assign rom[516][1] = -4;
assign rom[516][2] = 38;
assign rom[516][3] = -28;
assign rom[516][4] = -14;
assign rom[516][5] = 16;
assign rom[516][6] = -15;
assign rom[516][7] = -22;
assign rom[516][8] = -17;
assign rom[516][9] = -17;
assign rom[517][0] = -21;
assign rom[517][1] = 11;
assign rom[517][2] = 37;
assign rom[517][3] = -14;
assign rom[517][4] = -3;
assign rom[517][5] = 8;
assign rom[517][6] = -19;
assign rom[517][7] = -7;
assign rom[517][8] = -15;
assign rom[517][9] = -1;
assign rom[518][0] = -10;
assign rom[518][1] = 22;
assign rom[518][2] = 23;
assign rom[518][3] = -15;
assign rom[518][4] = 9;
assign rom[518][5] = 12;
assign rom[518][6] = -3;
assign rom[518][7] = 7;
assign rom[518][8] = -21;
assign rom[518][9] = -8;
assign rom[519][0] = -1;
assign rom[519][1] = 27;
assign rom[519][2] = -1;
assign rom[519][3] = -17;
assign rom[519][4] = 10;
assign rom[519][5] = 8;
assign rom[519][6] = 1;
assign rom[519][7] = 10;
assign rom[519][8] = -22;
assign rom[519][9] = 1;
assign rom[520][0] = -6;
assign rom[520][1] = 25;
assign rom[520][2] = -5;
assign rom[520][3] = 1;
assign rom[520][4] = -2;
assign rom[520][5] = 8;
assign rom[520][6] = -7;
assign rom[520][7] = 16;
assign rom[520][8] = -18;
assign rom[520][9] = -5;
assign rom[521][0] = -10;
assign rom[521][1] = 10;
assign rom[521][2] = 10;
assign rom[521][3] = 22;
assign rom[521][4] = 2;
assign rom[521][5] = -2;
assign rom[521][6] = -11;
assign rom[521][7] = -9;
assign rom[521][8] = -33;
assign rom[521][9] = -12;
assign rom[522][0] = -22;
assign rom[522][1] = 18;
assign rom[522][2] = 10;
assign rom[522][3] = 18;
assign rom[522][4] = -5;
assign rom[522][5] = 8;
assign rom[522][6] = -18;
assign rom[522][7] = -4;
assign rom[522][8] = -37;
assign rom[522][9] = -7;
assign rom[523][0] = -7;
assign rom[523][1] = 10;
assign rom[523][2] = 14;
assign rom[523][3] = 16;
assign rom[523][4] = -29;
assign rom[523][5] = -8;
assign rom[523][6] = -38;
assign rom[523][7] = -19;
assign rom[523][8] = -23;
assign rom[523][9] = -12;
assign rom[524][0] = 4;
assign rom[524][1] = 19;
assign rom[524][2] = 7;
assign rom[524][3] = 30;
assign rom[524][4] = -25;
assign rom[524][5] = -9;
assign rom[524][6] = -43;
assign rom[524][7] = -11;
assign rom[524][8] = -9;
assign rom[524][9] = -22;
assign rom[525][0] = 2;
assign rom[525][1] = 19;
assign rom[525][2] = 17;
assign rom[525][3] = 10;
assign rom[525][4] = -37;
assign rom[525][5] = 3;
assign rom[525][6] = -27;
assign rom[525][7] = -20;
assign rom[525][8] = 11;
assign rom[525][9] = -26;
assign rom[526][0] = 3;
assign rom[526][1] = 4;
assign rom[526][2] = 9;
assign rom[526][3] = 10;
assign rom[526][4] = -31;
assign rom[526][5] = 12;
assign rom[526][6] = -22;
assign rom[526][7] = -17;
assign rom[526][8] = 1;
assign rom[526][9] = -24;
assign rom[527][0] = 12;
assign rom[527][1] = 14;
assign rom[527][2] = 20;
assign rom[527][3] = 7;
assign rom[527][4] = -26;
assign rom[527][5] = 3;
assign rom[527][6] = -22;
assign rom[527][7] = -11;
assign rom[527][8] = 3;
assign rom[527][9] = -21;
assign rom[528][0] = 23;
assign rom[528][1] = 5;
assign rom[528][2] = 17;
assign rom[528][3] = 4;
assign rom[528][4] = -34;
assign rom[528][5] = 10;
assign rom[528][6] = -10;
assign rom[528][7] = -1;
assign rom[528][8] = -5;
assign rom[528][9] = -18;
assign rom[529][0] = 23;
assign rom[529][1] = -17;
assign rom[529][2] = 9;
assign rom[529][3] = -1;
assign rom[529][4] = -28;
assign rom[529][5] = 18;
assign rom[529][6] = -1;
assign rom[529][7] = -12;
assign rom[529][8] = -11;
assign rom[529][9] = -27;
assign rom[530][0] = 22;
assign rom[530][1] = -27;
assign rom[530][2] = 8;
assign rom[530][3] = 0;
assign rom[530][4] = -20;
assign rom[530][5] = 16;
assign rom[530][6] = 12;
assign rom[530][7] = 7;
assign rom[530][8] = 3;
assign rom[530][9] = -17;
assign rom[531][0] = 21;
assign rom[531][1] = -29;
assign rom[531][2] = 5;
assign rom[531][3] = 1;
assign rom[531][4] = -12;
assign rom[531][5] = -1;
assign rom[531][6] = 25;
assign rom[531][7] = -3;
assign rom[531][8] = 7;
assign rom[531][9] = -18;
assign rom[532][0] = 6;
assign rom[532][1] = -21;
assign rom[532][2] = -2;
assign rom[532][3] = -10;
assign rom[532][4] = -16;
assign rom[532][5] = 2;
assign rom[532][6] = 17;
assign rom[532][7] = -1;
assign rom[532][8] = 7;
assign rom[532][9] = -7;
assign rom[533][0] = 9;
assign rom[533][1] = -14;
assign rom[533][2] = -13;
assign rom[533][3] = 0;
assign rom[533][4] = -14;
assign rom[533][5] = 5;
assign rom[533][6] = 20;
assign rom[533][7] = -5;
assign rom[533][8] = -1;
assign rom[533][9] = -19;
assign rom[534][0] = 16;
assign rom[534][1] = -1;
assign rom[534][2] = -7;
assign rom[534][3] = 13;
assign rom[534][4] = 0;
assign rom[534][5] = 11;
assign rom[534][6] = 21;
assign rom[534][7] = -4;
assign rom[534][8] = -6;
assign rom[534][9] = -21;
assign rom[535][0] = 9;
assign rom[535][1] = 15;
assign rom[535][2] = 4;
assign rom[535][3] = 5;
assign rom[535][4] = -2;
assign rom[535][5] = 13;
assign rom[535][6] = 3;
assign rom[535][7] = -21;
assign rom[535][8] = -1;
assign rom[535][9] = -8;
assign rom[536][0] = -12;
assign rom[536][1] = 19;
assign rom[536][2] = 10;
assign rom[536][3] = 6;
assign rom[536][4] = 6;
assign rom[536][5] = 12;
assign rom[536][6] = 6;
assign rom[536][7] = -21;
assign rom[536][8] = 1;
assign rom[536][9] = -26;
assign rom[537][0] = -6;
assign rom[537][1] = 4;
assign rom[537][2] = 21;
assign rom[537][3] = 8;
assign rom[537][4] = -2;
assign rom[537][5] = 4;
assign rom[537][6] = 8;
assign rom[537][7] = -33;
assign rom[537][8] = -5;
assign rom[537][9] = -11;
assign rom[538][0] = 2;
assign rom[538][1] = -3;
assign rom[538][2] = 20;
assign rom[538][3] = 16;
assign rom[538][4] = -8;
assign rom[538][5] = 11;
assign rom[538][6] = -1;
assign rom[538][7] = -33;
assign rom[538][8] = -5;
assign rom[538][9] = -3;
assign rom[539][0] = -5;
assign rom[539][1] = -16;
assign rom[539][2] = 14;
assign rom[539][3] = -1;
assign rom[539][4] = 4;
assign rom[539][5] = 6;
assign rom[539][6] = -4;
assign rom[539][7] = -49;
assign rom[539][8] = 1;
assign rom[539][9] = -5;
assign rom[540][0] = -2;
assign rom[540][1] = -30;
assign rom[540][2] = 20;
assign rom[540][3] = -1;
assign rom[540][4] = -11;
assign rom[540][5] = 11;
assign rom[540][6] = -18;
assign rom[540][7] = -41;
assign rom[540][8] = -3;
assign rom[540][9] = -2;
assign rom[541][0] = -12;
assign rom[541][1] = -20;
assign rom[541][2] = 36;
assign rom[541][3] = -26;
assign rom[541][4] = -4;
assign rom[541][5] = 4;
assign rom[541][6] = -27;
assign rom[541][7] = -36;
assign rom[541][8] = -7;
assign rom[541][9] = 3;
assign rom[542][0] = -19;
assign rom[542][1] = -3;
assign rom[542][2] = 30;
assign rom[542][3] = -23;
assign rom[542][4] = -2;
assign rom[542][5] = 13;
assign rom[542][6] = -22;
assign rom[542][7] = -22;
assign rom[542][8] = -9;
assign rom[542][9] = 2;
assign rom[543][0] = -13;
assign rom[543][1] = 11;
assign rom[543][2] = 28;
assign rom[543][3] = -20;
assign rom[543][4] = -8;
assign rom[543][5] = 10;
assign rom[543][6] = -8;
assign rom[543][7] = -5;
assign rom[543][8] = -21;
assign rom[543][9] = 6;
assign rom[544][0] = -8;
assign rom[544][1] = 26;
assign rom[544][2] = 5;
assign rom[544][3] = -22;
assign rom[544][4] = 8;
assign rom[544][5] = 7;
assign rom[544][6] = -13;
assign rom[544][7] = 9;
assign rom[544][8] = -23;
assign rom[544][9] = -10;
assign rom[545][0] = -6;
assign rom[545][1] = 21;
assign rom[545][2] = 4;
assign rom[545][3] = -13;
assign rom[545][4] = 7;
assign rom[545][5] = 9;
assign rom[545][6] = 4;
assign rom[545][7] = 13;
assign rom[545][8] = -19;
assign rom[545][9] = -7;
assign rom[546][0] = -8;
assign rom[546][1] = 28;
assign rom[546][2] = -2;
assign rom[546][3] = -3;
assign rom[546][4] = 3;
assign rom[546][5] = 20;
assign rom[546][6] = -7;
assign rom[546][7] = 8;
assign rom[546][8] = -25;
assign rom[546][9] = -9;
assign rom[547][0] = -13;
assign rom[547][1] = 11;
assign rom[547][2] = -1;
assign rom[547][3] = 8;
assign rom[547][4] = 5;
assign rom[547][5] = 1;
assign rom[547][6] = -3;
assign rom[547][7] = -6;
assign rom[547][8] = -19;
assign rom[547][9] = -14;
assign rom[548][0] = -19;
assign rom[548][1] = 16;
assign rom[548][2] = -1;
assign rom[548][3] = 18;
assign rom[548][4] = -11;
assign rom[548][5] = 6;
assign rom[548][6] = -16;
assign rom[548][7] = -10;
assign rom[548][8] = -39;
assign rom[548][9] = -13;
assign rom[549][0] = -16;
assign rom[549][1] = 26;
assign rom[549][2] = 12;
assign rom[549][3] = 15;
assign rom[549][4] = -26;
assign rom[549][5] = 1;
assign rom[549][6] = -29;
assign rom[549][7] = 6;
assign rom[549][8] = -34;
assign rom[549][9] = -19;
assign rom[550][0] = -4;
assign rom[550][1] = 21;
assign rom[550][2] = 11;
assign rom[550][3] = 25;
assign rom[550][4] = -18;
assign rom[550][5] = -10;
assign rom[550][6] = -38;
assign rom[550][7] = 7;
assign rom[550][8] = -14;
assign rom[550][9] = -28;
assign rom[551][0] = -5;
assign rom[551][1] = 19;
assign rom[551][2] = 11;
assign rom[551][3] = 14;
assign rom[551][4] = -24;
assign rom[551][5] = -11;
assign rom[551][6] = -37;
assign rom[551][7] = 5;
assign rom[551][8] = -10;
assign rom[551][9] = -21;
assign rom[552][0] = 7;
assign rom[552][1] = 16;
assign rom[552][2] = -1;
assign rom[552][3] = 10;
assign rom[552][4] = -24;
assign rom[552][5] = 3;
assign rom[552][6] = -23;
assign rom[552][7] = 6;
assign rom[552][8] = 4;
assign rom[552][9] = -20;
assign rom[553][0] = 13;
assign rom[553][1] = 4;
assign rom[553][2] = 9;
assign rom[553][3] = 15;
assign rom[553][4] = -23;
assign rom[553][5] = 0;
assign rom[553][6] = -22;
assign rom[553][7] = -10;
assign rom[553][8] = -5;
assign rom[553][9] = -22;
assign rom[554][0] = 12;
assign rom[554][1] = 1;
assign rom[554][2] = 11;
assign rom[554][3] = 12;
assign rom[554][4] = -15;
assign rom[554][5] = 3;
assign rom[554][6] = -17;
assign rom[554][7] = -1;
assign rom[554][8] = 3;
assign rom[554][9] = -18;
assign rom[555][0] = 24;
assign rom[555][1] = -3;
assign rom[555][2] = 6;
assign rom[555][3] = 2;
assign rom[555][4] = -1;
assign rom[555][5] = 7;
assign rom[555][6] = -18;
assign rom[555][7] = -9;
assign rom[555][8] = 3;
assign rom[555][9] = -7;
assign rom[556][0] = 23;
assign rom[556][1] = -17;
assign rom[556][2] = 2;
assign rom[556][3] = 8;
assign rom[556][4] = -10;
assign rom[556][5] = 7;
assign rom[556][6] = -13;
assign rom[556][7] = -10;
assign rom[556][8] = 24;
assign rom[556][9] = -14;
assign rom[557][0] = 26;
assign rom[557][1] = -31;
assign rom[557][2] = 0;
assign rom[557][3] = 3;
assign rom[557][4] = -12;
assign rom[557][5] = 8;
assign rom[557][6] = -8;
assign rom[557][7] = -8;
assign rom[557][8] = 21;
assign rom[557][9] = -14;
assign rom[558][0] = 24;
assign rom[558][1] = -9;
assign rom[558][2] = -14;
assign rom[558][3] = -9;
assign rom[558][4] = -9;
assign rom[558][5] = 17;
assign rom[558][6] = 0;
assign rom[558][7] = -5;
assign rom[558][8] = 22;
assign rom[558][9] = -19;
assign rom[559][0] = 16;
assign rom[559][1] = 6;
assign rom[559][2] = -16;
assign rom[559][3] = -1;
assign rom[559][4] = -4;
assign rom[559][5] = 15;
assign rom[559][6] = -7;
assign rom[559][7] = 0;
assign rom[559][8] = 12;
assign rom[559][9] = -23;
assign rom[560][0] = 6;
assign rom[560][1] = 15;
assign rom[560][2] = -2;
assign rom[560][3] = 3;
assign rom[560][4] = -5;
assign rom[560][5] = 4;
assign rom[560][6] = 1;
assign rom[560][7] = 3;
assign rom[560][8] = 12;
assign rom[560][9] = -19;
assign rom[561][0] = 12;
assign rom[561][1] = 12;
assign rom[561][2] = 6;
assign rom[561][3] = 10;
assign rom[561][4] = 1;
assign rom[561][5] = -5;
assign rom[561][6] = -2;
assign rom[561][7] = -9;
assign rom[561][8] = 12;
assign rom[561][9] = -11;
assign rom[562][0] = 0;
assign rom[562][1] = 24;
assign rom[562][2] = -2;
assign rom[562][3] = 0;
assign rom[562][4] = 14;
assign rom[562][5] = 2;
assign rom[562][6] = -12;
assign rom[562][7] = -7;
assign rom[562][8] = 3;
assign rom[562][9] = -21;
assign rom[563][0] = -18;
assign rom[563][1] = 3;
assign rom[563][2] = 7;
assign rom[563][3] = 5;
assign rom[563][4] = 21;
assign rom[563][5] = 5;
assign rom[563][6] = -10;
assign rom[563][7] = -25;
assign rom[563][8] = -3;
assign rom[563][9] = -24;
assign rom[564][0] = -20;
assign rom[564][1] = -13;
assign rom[564][2] = 7;
assign rom[564][3] = -2;
assign rom[564][4] = 14;
assign rom[564][5] = 8;
assign rom[564][6] = -20;
assign rom[564][7] = -34;
assign rom[564][8] = 8;
assign rom[564][9] = -15;
assign rom[565][0] = -18;
assign rom[565][1] = -12;
assign rom[565][2] = 20;
assign rom[565][3] = -4;
assign rom[565][4] = 14;
assign rom[565][5] = 12;
assign rom[565][6] = -16;
assign rom[565][7] = -43;
assign rom[565][8] = -1;
assign rom[565][9] = -4;
assign rom[566][0] = -23;
assign rom[566][1] = -6;
assign rom[566][2] = 26;
assign rom[566][3] = -24;
assign rom[566][4] = 7;
assign rom[566][5] = 11;
assign rom[566][6] = -23;
assign rom[566][7] = -29;
assign rom[566][8] = -1;
assign rom[566][9] = 17;
assign rom[567][0] = -21;
assign rom[567][1] = -6;
assign rom[567][2] = 19;
assign rom[567][3] = -17;
assign rom[567][4] = -1;
assign rom[567][5] = 15;
assign rom[567][6] = -23;
assign rom[567][7] = -18;
assign rom[567][8] = -3;
assign rom[567][9] = 6;
assign rom[568][0] = -16;
assign rom[568][1] = 12;
assign rom[568][2] = 17;
assign rom[568][3] = -18;
assign rom[568][4] = 7;
assign rom[568][5] = 21;
assign rom[568][6] = -15;
assign rom[568][7] = -13;
assign rom[568][8] = -20;
assign rom[568][9] = 1;
assign rom[569][0] = -12;
assign rom[569][1] = 7;
assign rom[569][2] = 14;
assign rom[569][3] = -13;
assign rom[569][4] = -1;
assign rom[569][5] = 23;
assign rom[569][6] = -3;
assign rom[569][7] = 7;
assign rom[569][8] = -21;
assign rom[569][9] = 1;
assign rom[570][0] = -17;
assign rom[570][1] = 16;
assign rom[570][2] = 8;
assign rom[570][3] = -7;
assign rom[570][4] = 7;
assign rom[570][5] = 20;
assign rom[570][6] = -12;
assign rom[570][7] = 2;
assign rom[570][8] = -22;
assign rom[570][9] = 2;
assign rom[571][0] = -16;
assign rom[571][1] = 19;
assign rom[571][2] = -9;
assign rom[571][3] = -16;
assign rom[571][4] = 4;
assign rom[571][5] = 11;
assign rom[571][6] = -5;
assign rom[571][7] = 18;
assign rom[571][8] = -31;
assign rom[571][9] = -10;
assign rom[572][0] = -3;
assign rom[572][1] = 26;
assign rom[572][2] = -8;
assign rom[572][3] = -15;
assign rom[572][4] = 14;
assign rom[572][5] = 22;
assign rom[572][6] = -3;
assign rom[572][7] = 3;
assign rom[572][8] = -28;
assign rom[572][9] = 6;
assign rom[573][0] = -1;
assign rom[573][1] = 13;
assign rom[573][2] = -15;
assign rom[573][3] = 10;
assign rom[573][4] = 10;
assign rom[573][5] = 17;
assign rom[573][6] = -6;
assign rom[573][7] = -1;
assign rom[573][8] = -21;
assign rom[573][9] = -12;
assign rom[574][0] = -20;
assign rom[574][1] = 20;
assign rom[574][2] = -6;
assign rom[574][3] = 24;
assign rom[574][4] = -8;
assign rom[574][5] = 2;
assign rom[574][6] = -12;
assign rom[574][7] = -2;
assign rom[574][8] = -39;
assign rom[574][9] = -20;
assign rom[575][0] = -17;
assign rom[575][1] = 12;
assign rom[575][2] = -15;
assign rom[575][3] = 19;
assign rom[575][4] = -8;
assign rom[575][5] = 8;
assign rom[575][6] = -3;
assign rom[575][7] = 22;
assign rom[575][8] = -44;
assign rom[575][9] = -17;
assign rom[576][0] = -20;
assign rom[576][1] = 15;
assign rom[576][2] = -18;
assign rom[576][3] = 18;
assign rom[576][4] = -13;
assign rom[576][5] = -10;
assign rom[576][6] = -15;
assign rom[576][7] = 24;
assign rom[576][8] = -24;
assign rom[576][9] = -8;
assign rom[577][0] = 1;
assign rom[577][1] = 8;
assign rom[577][2] = -5;
assign rom[577][3] = 22;
assign rom[577][4] = -11;
assign rom[577][5] = -12;
assign rom[577][6] = -31;
assign rom[577][7] = 17;
assign rom[577][8] = -22;
assign rom[577][9] = -7;
assign rom[578][0] = 5;
assign rom[578][1] = -2;
assign rom[578][2] = -17;
assign rom[578][3] = 11;
assign rom[578][4] = -15;
assign rom[578][5] = -2;
assign rom[578][6] = -29;
assign rom[578][7] = 17;
assign rom[578][8] = -7;
assign rom[578][9] = -3;
assign rom[579][0] = 2;
assign rom[579][1] = 6;
assign rom[579][2] = -4;
assign rom[579][3] = 12;
assign rom[579][4] = -14;
assign rom[579][5] = -6;
assign rom[579][6] = -33;
assign rom[579][7] = 19;
assign rom[579][8] = 6;
assign rom[579][9] = 2;
assign rom[580][0] = 1;
assign rom[580][1] = -3;
assign rom[580][2] = -4;
assign rom[580][3] = 6;
assign rom[580][4] = 2;
assign rom[580][5] = 3;
assign rom[580][6] = -22;
assign rom[580][7] = -3;
assign rom[580][8] = 6;
assign rom[580][9] = -6;
assign rom[581][0] = 20;
assign rom[581][1] = -23;
assign rom[581][2] = 0;
assign rom[581][3] = 4;
assign rom[581][4] = -2;
assign rom[581][5] = 8;
assign rom[581][6] = -21;
assign rom[581][7] = 1;
assign rom[581][8] = 5;
assign rom[581][9] = -15;
assign rom[582][0] = 13;
assign rom[582][1] = -20;
assign rom[582][2] = -1;
assign rom[582][3] = 8;
assign rom[582][4] = -2;
assign rom[582][5] = 14;
assign rom[582][6] = -31;
assign rom[582][7] = -5;
assign rom[582][8] = 11;
assign rom[582][9] = -7;
assign rom[583][0] = 23;
assign rom[583][1] = -23;
assign rom[583][2] = -9;
assign rom[583][3] = 1;
assign rom[583][4] = -15;
assign rom[583][5] = 20;
assign rom[583][6] = -27;
assign rom[583][7] = 3;
assign rom[583][8] = 18;
assign rom[583][9] = -8;
assign rom[584][0] = 15;
assign rom[584][1] = -24;
assign rom[584][2] = -4;
assign rom[584][3] = 10;
assign rom[584][4] = -8;
assign rom[584][5] = 2;
assign rom[584][6] = -32;
assign rom[584][7] = 7;
assign rom[584][8] = 27;
assign rom[584][9] = -14;
assign rom[585][0] = 19;
assign rom[585][1] = -13;
assign rom[585][2] = -8;
assign rom[585][3] = -2;
assign rom[585][4] = 5;
assign rom[585][5] = 14;
assign rom[585][6] = -21;
assign rom[585][7] = 0;
assign rom[585][8] = 13;
assign rom[585][9] = -14;
assign rom[586][0] = 4;
assign rom[586][1] = 3;
assign rom[586][2] = -14;
assign rom[586][3] = -3;
assign rom[586][4] = 4;
assign rom[586][5] = 1;
assign rom[586][6] = -18;
assign rom[586][7] = 11;
assign rom[586][8] = 22;
assign rom[586][9] = -7;
assign rom[587][0] = -4;
assign rom[587][1] = 24;
assign rom[587][2] = -17;
assign rom[587][3] = 0;
assign rom[587][4] = 0;
assign rom[587][5] = 0;
assign rom[587][6] = -27;
assign rom[587][7] = 1;
assign rom[587][8] = 5;
assign rom[587][9] = -14;
assign rom[588][0] = -16;
assign rom[588][1] = 27;
assign rom[588][2] = -4;
assign rom[588][3] = -1;
assign rom[588][4] = 5;
assign rom[588][5] = -12;
assign rom[588][6] = -31;
assign rom[588][7] = -6;
assign rom[588][8] = 14;
assign rom[588][9] = 1;
assign rom[589][0] = -19;
assign rom[589][1] = 19;
assign rom[589][2] = 1;
assign rom[589][3] = -2;
assign rom[589][4] = 12;
assign rom[589][5] = -7;
assign rom[589][6] = -16;
assign rom[589][7] = -13;
assign rom[589][8] = 14;
assign rom[589][9] = 6;
assign rom[590][0] = -25;
assign rom[590][1] = 6;
assign rom[590][2] = -2;
assign rom[590][3] = -11;
assign rom[590][4] = 16;
assign rom[590][5] = -4;
assign rom[590][6] = -27;
assign rom[590][7] = -26;
assign rom[590][8] = 15;
assign rom[590][9] = 13;
assign rom[591][0] = -30;
assign rom[591][1] = -11;
assign rom[591][2] = 6;
assign rom[591][3] = -7;
assign rom[591][4] = 17;
assign rom[591][5] = 7;
assign rom[591][6] = -24;
assign rom[591][7] = -34;
assign rom[591][8] = 7;
assign rom[591][9] = 24;
assign rom[592][0] = -17;
assign rom[592][1] = -4;
assign rom[592][2] = 5;
assign rom[592][3] = -29;
assign rom[592][4] = 17;
assign rom[592][5] = -5;
assign rom[592][6] = -21;
assign rom[592][7] = -23;
assign rom[592][8] = -12;
assign rom[592][9] = 23;
assign rom[593][0] = -10;
assign rom[593][1] = 4;
assign rom[593][2] = 13;
assign rom[593][3] = -27;
assign rom[593][4] = -6;
assign rom[593][5] = 0;
assign rom[593][6] = -9;
assign rom[593][7] = -22;
assign rom[593][8] = -10;
assign rom[593][9] = 11;
assign rom[594][0] = -8;
assign rom[594][1] = 18;
assign rom[594][2] = 3;
assign rom[594][3] = -12;
assign rom[594][4] = 7;
assign rom[594][5] = 15;
assign rom[594][6] = -21;
assign rom[594][7] = -19;
assign rom[594][8] = -14;
assign rom[594][9] = 10;
assign rom[595][0] = -16;
assign rom[595][1] = 15;
assign rom[595][2] = 3;
assign rom[595][3] = -22;
assign rom[595][4] = -1;
assign rom[595][5] = 16;
assign rom[595][6] = -10;
assign rom[595][7] = 6;
assign rom[595][8] = -20;
assign rom[595][9] = 5;
assign rom[596][0] = -13;
assign rom[596][1] = 29;
assign rom[596][2] = -6;
assign rom[596][3] = -6;
assign rom[596][4] = 15;
assign rom[596][5] = 18;
assign rom[596][6] = -1;
assign rom[596][7] = 11;
assign rom[596][8] = -33;
assign rom[596][9] = -3;
assign rom[597][0] = -11;
assign rom[597][1] = 18;
assign rom[597][2] = 5;
assign rom[597][3] = -21;
assign rom[597][4] = 13;
assign rom[597][5] = 15;
assign rom[597][6] = -10;
assign rom[597][7] = 5;
assign rom[597][8] = -21;
assign rom[597][9] = -7;
assign rom[598][0] = -12;
assign rom[598][1] = 21;
assign rom[598][2] = 6;
assign rom[598][3] = -8;
assign rom[598][4] = 14;
assign rom[598][5] = 17;
assign rom[598][6] = -8;
assign rom[598][7] = 18;
assign rom[598][8] = -29;
assign rom[598][9] = -5;
assign rom[599][0] = -12;
assign rom[599][1] = 17;
assign rom[599][2] = -14;
assign rom[599][3] = -9;
assign rom[599][4] = 4;
assign rom[599][5] = 14;
assign rom[599][6] = -8;
assign rom[599][7] = 17;
assign rom[599][8] = -16;
assign rom[599][9] = -11;
assign rom[600][0] = -10;
assign rom[600][1] = 17;
assign rom[600][2] = -9;
assign rom[600][3] = 6;
assign rom[600][4] = 6;
assign rom[600][5] = 11;
assign rom[600][6] = 6;
assign rom[600][7] = 11;
assign rom[600][8] = -24;
assign rom[600][9] = 4;
assign rom[601][0] = -19;
assign rom[601][1] = 13;
assign rom[601][2] = -17;
assign rom[601][3] = 24;
assign rom[601][4] = -4;
assign rom[601][5] = 9;
assign rom[601][6] = -3;
assign rom[601][7] = 19;
assign rom[601][8] = -30;
assign rom[601][9] = -1;
assign rom[602][0] = -26;
assign rom[602][1] = 13;
assign rom[602][2] = -33;
assign rom[602][3] = 29;
assign rom[602][4] = -11;
assign rom[602][5] = -10;
assign rom[602][6] = -8;
assign rom[602][7] = 26;
assign rom[602][8] = -51;
assign rom[602][9] = -1;
assign rom[603][0] = -17;
assign rom[603][1] = -2;
assign rom[603][2] = -33;
assign rom[603][3] = 20;
assign rom[603][4] = -13;
assign rom[603][5] = -3;
assign rom[603][6] = -14;
assign rom[603][7] = 31;
assign rom[603][8] = -42;
assign rom[603][9] = 18;
assign rom[604][0] = -27;
assign rom[604][1] = -22;
assign rom[604][2] = -30;
assign rom[604][3] = 23;
assign rom[604][4] = -16;
assign rom[604][5] = -4;
assign rom[604][6] = -23;
assign rom[604][7] = 32;
assign rom[604][8] = -19;
assign rom[604][9] = 6;
assign rom[605][0] = -21;
assign rom[605][1] = -13;
assign rom[605][2] = -29;
assign rom[605][3] = 21;
assign rom[605][4] = -15;
assign rom[605][5] = -2;
assign rom[605][6] = -23;
assign rom[605][7] = 11;
assign rom[605][8] = -18;
assign rom[605][9] = 15;
assign rom[606][0] = -18;
assign rom[606][1] = -32;
assign rom[606][2] = -19;
assign rom[606][3] = 15;
assign rom[606][4] = -23;
assign rom[606][5] = 0;
assign rom[606][6] = -24;
assign rom[606][7] = 11;
assign rom[606][8] = -10;
assign rom[606][9] = 3;
assign rom[607][0] = -12;
assign rom[607][1] = -29;
assign rom[607][2] = -20;
assign rom[607][3] = 19;
assign rom[607][4] = -15;
assign rom[607][5] = 2;
assign rom[607][6] = -41;
assign rom[607][7] = 18;
assign rom[607][8] = -9;
assign rom[607][9] = 15;
assign rom[608][0] = -8;
assign rom[608][1] = -37;
assign rom[608][2] = -18;
assign rom[608][3] = 18;
assign rom[608][4] = -14;
assign rom[608][5] = 7;
assign rom[608][6] = -28;
assign rom[608][7] = 20;
assign rom[608][8] = 2;
assign rom[608][9] = 0;
assign rom[609][0] = -4;
assign rom[609][1] = -41;
assign rom[609][2] = -3;
assign rom[609][3] = 13;
assign rom[609][4] = -23;
assign rom[609][5] = 8;
assign rom[609][6] = -27;
assign rom[609][7] = 9;
assign rom[609][8] = 10;
assign rom[609][9] = 4;
assign rom[610][0] = -7;
assign rom[610][1] = -32;
assign rom[610][2] = -18;
assign rom[610][3] = 8;
assign rom[610][4] = -18;
assign rom[610][5] = 13;
assign rom[610][6] = -37;
assign rom[610][7] = 21;
assign rom[610][8] = 12;
assign rom[610][9] = 1;
assign rom[611][0] = -5;
assign rom[611][1] = -37;
assign rom[611][2] = -10;
assign rom[611][3] = 9;
assign rom[611][4] = -23;
assign rom[611][5] = 8;
assign rom[611][6] = -33;
assign rom[611][7] = 19;
assign rom[611][8] = 14;
assign rom[611][9] = -5;
assign rom[612][0] = -17;
assign rom[612][1] = -24;
assign rom[612][2] = -22;
assign rom[612][3] = 13;
assign rom[612][4] = -12;
assign rom[612][5] = 0;
assign rom[612][6] = -29;
assign rom[612][7] = 26;
assign rom[612][8] = 13;
assign rom[612][9] = -5;
assign rom[613][0] = -19;
assign rom[613][1] = 2;
assign rom[613][2] = -21;
assign rom[613][3] = 4;
assign rom[613][4] = -29;
assign rom[613][5] = 5;
assign rom[613][6] = -30;
assign rom[613][7] = 8;
assign rom[613][8] = 12;
assign rom[613][9] = 3;
assign rom[614][0] = -24;
assign rom[614][1] = 11;
assign rom[614][2] = -6;
assign rom[614][3] = -9;
assign rom[614][4] = -21;
assign rom[614][5] = -1;
assign rom[614][6] = -33;
assign rom[614][7] = 5;
assign rom[614][8] = 8;
assign rom[614][9] = 13;
assign rom[615][0] = -22;
assign rom[615][1] = 21;
assign rom[615][2] = -19;
assign rom[615][3] = -13;
assign rom[615][4] = -18;
assign rom[615][5] = -8;
assign rom[615][6] = -25;
assign rom[615][7] = -8;
assign rom[615][8] = 17;
assign rom[615][9] = 8;
assign rom[616][0] = -37;
assign rom[616][1] = 18;
assign rom[616][2] = -3;
assign rom[616][3] = -15;
assign rom[616][4] = 3;
assign rom[616][5] = -16;
assign rom[616][6] = -24;
assign rom[616][7] = -11;
assign rom[616][8] = 12;
assign rom[616][9] = 29;
assign rom[617][0] = -27;
assign rom[617][1] = 19;
assign rom[617][2] = -11;
assign rom[617][3] = -21;
assign rom[617][4] = -12;
assign rom[617][5] = 4;
assign rom[617][6] = -11;
assign rom[617][7] = -5;
assign rom[617][8] = 5;
assign rom[617][9] = 21;
assign rom[618][0] = -23;
assign rom[618][1] = 9;
assign rom[618][2] = -4;
assign rom[618][3] = -16;
assign rom[618][4] = 9;
assign rom[618][5] = 10;
assign rom[618][6] = -24;
assign rom[618][7] = -21;
assign rom[618][8] = -13;
assign rom[618][9] = 25;
assign rom[619][0] = -21;
assign rom[619][1] = 8;
assign rom[619][2] = -10;
assign rom[619][3] = -16;
assign rom[619][4] = -5;
assign rom[619][5] = 18;
assign rom[619][6] = -15;
assign rom[619][7] = -13;
assign rom[619][8] = -16;
assign rom[619][9] = 19;
assign rom[620][0] = -10;
assign rom[620][1] = 24;
assign rom[620][2] = 0;
assign rom[620][3] = -16;
assign rom[620][4] = -5;
assign rom[620][5] = 16;
assign rom[620][6] = 0;
assign rom[620][7] = -1;
assign rom[620][8] = -17;
assign rom[620][9] = 19;
assign rom[621][0] = -16;
assign rom[621][1] = 25;
assign rom[621][2] = 4;
assign rom[621][3] = -21;
assign rom[621][4] = 9;
assign rom[621][5] = 11;
assign rom[621][6] = 4;
assign rom[621][7] = 8;
assign rom[621][8] = -30;
assign rom[621][9] = -6;
assign rom[622][0] = -1;
assign rom[622][1] = 28;
assign rom[622][2] = 4;
assign rom[622][3] = -18;
assign rom[622][4] = 5;
assign rom[622][5] = 16;
assign rom[622][6] = -3;
assign rom[622][7] = 10;
assign rom[622][8] = -26;
assign rom[622][9] = -6;
assign rom[623][0] = 1;
assign rom[623][1] = 32;
assign rom[623][2] = -9;
assign rom[623][3] = -14;
assign rom[623][4] = 5;
assign rom[623][5] = 9;
assign rom[623][6] = 5;
assign rom[623][7] = 6;
assign rom[623][8] = -21;
assign rom[623][9] = -4;
assign rom[624][0] = -8;
assign rom[624][1] = 29;
assign rom[624][2] = -9;
assign rom[624][3] = -20;
assign rom[624][4] = 9;
assign rom[624][5] = 17;
assign rom[624][6] = 0;
assign rom[624][7] = 20;
assign rom[624][8] = -17;
assign rom[624][9] = -4;
assign rom[625][0] = -15;
assign rom[625][1] = 32;
assign rom[625][2] = -12;
assign rom[625][3] = -17;
assign rom[625][4] = 2;
assign rom[625][5] = 17;
assign rom[625][6] = -3;
assign rom[625][7] = 13;
assign rom[625][8] = -27;
assign rom[625][9] = 0;
assign rom[626][0] = -15;
assign rom[626][1] = 15;
assign rom[626][2] = -2;
assign rom[626][3] = -15;
assign rom[626][4] = 0;
assign rom[626][5] = 18;
assign rom[626][6] = -9;
assign rom[626][7] = 13;
assign rom[626][8] = -22;
assign rom[626][9] = 0;
assign rom[627][0] = -6;
assign rom[627][1] = 16;
assign rom[627][2] = -12;
assign rom[627][3] = -6;
assign rom[627][4] = -6;
assign rom[627][5] = 20;
assign rom[627][6] = 6;
assign rom[627][7] = 12;
assign rom[627][8] = -39;
assign rom[627][9] = 7;
assign rom[628][0] = -17;
assign rom[628][1] = 2;
assign rom[628][2] = -20;
assign rom[628][3] = 2;
assign rom[628][4] = -8;
assign rom[628][5] = -4;
assign rom[628][6] = -7;
assign rom[628][7] = 22;
assign rom[628][8] = -36;
assign rom[628][9] = 11;
assign rom[629][0] = -30;
assign rom[629][1] = -6;
assign rom[629][2] = -35;
assign rom[629][3] = 23;
assign rom[629][4] = -26;
assign rom[629][5] = 3;
assign rom[629][6] = -7;
assign rom[629][7] = 16;
assign rom[629][8] = -40;
assign rom[629][9] = 17;
assign rom[630][0] = -34;
assign rom[630][1] = -5;
assign rom[630][2] = -38;
assign rom[630][3] = 13;
assign rom[630][4] = -20;
assign rom[630][5] = -15;
assign rom[630][6] = -12;
assign rom[630][7] = 23;
assign rom[630][8] = -33;
assign rom[630][9] = 19;
assign rom[631][0] = -35;
assign rom[631][1] = -15;
assign rom[631][2] = -25;
assign rom[631][3] = 16;
assign rom[631][4] = -28;
assign rom[631][5] = -14;
assign rom[631][6] = -20;
assign rom[631][7] = 25;
assign rom[631][8] = -31;
assign rom[631][9] = 5;
assign rom[632][0] = -46;
assign rom[632][1] = -26;
assign rom[632][2] = -37;
assign rom[632][3] = 22;
assign rom[632][4] = -34;
assign rom[632][5] = -1;
assign rom[632][6] = -10;
assign rom[632][7] = 15;
assign rom[632][8] = -38;
assign rom[632][9] = 20;
assign rom[633][0] = -33;
assign rom[633][1] = -33;
assign rom[633][2] = -26;
assign rom[633][3] = 33;
assign rom[633][4] = -37;
assign rom[633][5] = 8;
assign rom[633][6] = -21;
assign rom[633][7] = 26;
assign rom[633][8] = -26;
assign rom[633][9] = 20;
assign rom[634][0] = -32;
assign rom[634][1] = -38;
assign rom[634][2] = -30;
assign rom[634][3] = 23;
assign rom[634][4] = -43;
assign rom[634][5] = 10;
assign rom[634][6] = -15;
assign rom[634][7] = 19;
assign rom[634][8] = -26;
assign rom[634][9] = 24;
assign rom[635][0] = -34;
assign rom[635][1] = -40;
assign rom[635][2] = -20;
assign rom[635][3] = 21;
assign rom[635][4] = -50;
assign rom[635][5] = 4;
assign rom[635][6] = -16;
assign rom[635][7] = 14;
assign rom[635][8] = -35;
assign rom[635][9] = 13;
assign rom[636][0] = -34;
assign rom[636][1] = -30;
assign rom[636][2] = -19;
assign rom[636][3] = 28;
assign rom[636][4] = -34;
assign rom[636][5] = 3;
assign rom[636][6] = -31;
assign rom[636][7] = 15;
assign rom[636][8] = -19;
assign rom[636][9] = 17;
assign rom[637][0] = -33;
assign rom[637][1] = -37;
assign rom[637][2] = -21;
assign rom[637][3] = 10;
assign rom[637][4] = -37;
assign rom[637][5] = 4;
assign rom[637][6] = -27;
assign rom[637][7] = 20;
assign rom[637][8] = -14;
assign rom[637][9] = 4;
assign rom[638][0] = -38;
assign rom[638][1] = -21;
assign rom[638][2] = -20;
assign rom[638][3] = 6;
assign rom[638][4] = -50;
assign rom[638][5] = 2;
assign rom[638][6] = -23;
assign rom[638][7] = 20;
assign rom[638][8] = -16;
assign rom[638][9] = 10;
assign rom[639][0] = -41;
assign rom[639][1] = -14;
assign rom[639][2] = -18;
assign rom[639][3] = -4;
assign rom[639][4] = -39;
assign rom[639][5] = 9;
assign rom[639][6] = -28;
assign rom[639][7] = 19;
assign rom[639][8] = -2;
assign rom[639][9] = 30;
assign rom[640][0] = -24;
assign rom[640][1] = 8;
assign rom[640][2] = -22;
assign rom[640][3] = -11;
assign rom[640][4] = -38;
assign rom[640][5] = 1;
assign rom[640][6] = -12;
assign rom[640][7] = 22;
assign rom[640][8] = -14;
assign rom[640][9] = 27;
assign rom[641][0] = -38;
assign rom[641][1] = 15;
assign rom[641][2] = -15;
assign rom[641][3] = -2;
assign rom[641][4] = -33;
assign rom[641][5] = -9;
assign rom[641][6] = -17;
assign rom[641][7] = 20;
assign rom[641][8] = -12;
assign rom[641][9] = 26;
assign rom[642][0] = -23;
assign rom[642][1] = 22;
assign rom[642][2] = -25;
assign rom[642][3] = -5;
assign rom[642][4] = -37;
assign rom[642][5] = -12;
assign rom[642][6] = -16;
assign rom[642][7] = -1;
assign rom[642][8] = -13;
assign rom[642][9] = 31;
assign rom[643][0] = -22;
assign rom[643][1] = 23;
assign rom[643][2] = -15;
assign rom[643][3] = -10;
assign rom[643][4] = -23;
assign rom[643][5] = 3;
assign rom[643][6] = -8;
assign rom[643][7] = -4;
assign rom[643][8] = -12;
assign rom[643][9] = 38;
assign rom[644][0] = -22;
assign rom[644][1] = 22;
assign rom[644][2] = -7;
assign rom[644][3] = -14;
assign rom[644][4] = -7;
assign rom[644][5] = 0;
assign rom[644][6] = 2;
assign rom[644][7] = -1;
assign rom[644][8] = -28;
assign rom[644][9] = 37;
assign rom[645][0] = -19;
assign rom[645][1] = 14;
assign rom[645][2] = -15;
assign rom[645][3] = -19;
assign rom[645][4] = -3;
assign rom[645][5] = 8;
assign rom[645][6] = 3;
assign rom[645][7] = 8;
assign rom[645][8] = -29;
assign rom[645][9] = 19;
assign rom[646][0] = -16;
assign rom[646][1] = 14;
assign rom[646][2] = -13;
assign rom[646][3] = -6;
assign rom[646][4] = 4;
assign rom[646][5] = 23;
assign rom[646][6] = 2;
assign rom[646][7] = 5;
assign rom[646][8] = -26;
assign rom[646][9] = 10;
assign rom[647][0] = -3;
assign rom[647][1] = 16;
assign rom[647][2] = 1;
assign rom[647][3] = -19;
assign rom[647][4] = 3;
assign rom[647][5] = 15;
assign rom[647][6] = 6;
assign rom[647][7] = 0;
assign rom[647][8] = -19;
assign rom[647][9] = -1;
assign rom[648][0] = 0;
assign rom[648][1] = 17;
assign rom[648][2] = 6;
assign rom[648][3] = -17;
assign rom[648][4] = 3;
assign rom[648][5] = 18;
assign rom[648][6] = 2;
assign rom[648][7] = 4;
assign rom[648][8] = -16;
assign rom[648][9] = 4;
assign rom[649][0] = -12;
assign rom[649][1] = 16;
assign rom[649][2] = -5;
assign rom[649][3] = -5;
assign rom[649][4] = -1;
assign rom[649][5] = 21;
assign rom[649][6] = 7;
assign rom[649][7] = 7;
assign rom[649][8] = -21;
assign rom[649][9] = -2;
assign rom[650][0] = -13;
assign rom[650][1] = 16;
assign rom[650][2] = -6;
assign rom[650][3] = -19;
assign rom[650][4] = 4;
assign rom[650][5] = 8;
assign rom[650][6] = -2;
assign rom[650][7] = 11;
assign rom[650][8] = -16;
assign rom[650][9] = 0;
assign rom[651][0] = 1;
assign rom[651][1] = 24;
assign rom[651][2] = -8;
assign rom[651][3] = -11;
assign rom[651][4] = 6;
assign rom[651][5] = 12;
assign rom[651][6] = -2;
assign rom[651][7] = 5;
assign rom[651][8] = -18;
assign rom[651][9] = -10;
assign rom[652][0] = -12;
assign rom[652][1] = 29;
assign rom[652][2] = 2;
assign rom[652][3] = -22;
assign rom[652][4] = 2;
assign rom[652][5] = 12;
assign rom[652][6] = 4;
assign rom[652][7] = 5;
assign rom[652][8] = -18;
assign rom[652][9] = -5;
assign rom[653][0] = -11;
assign rom[653][1] = 27;
assign rom[653][2] = -1;
assign rom[653][3] = -7;
assign rom[653][4] = 2;
assign rom[653][5] = 19;
assign rom[653][6] = 3;
assign rom[653][7] = 12;
assign rom[653][8] = -26;
assign rom[653][9] = -7;
assign rom[654][0] = -14;
assign rom[654][1] = 19;
assign rom[654][2] = -4;
assign rom[654][3] = -14;
assign rom[654][4] = 7;
assign rom[654][5] = 10;
assign rom[654][6] = -2;
assign rom[654][7] = 8;
assign rom[654][8] = -33;
assign rom[654][9] = 14;
assign rom[655][0] = -5;
assign rom[655][1] = 23;
assign rom[655][2] = -8;
assign rom[655][3] = -15;
assign rom[655][4] = 3;
assign rom[655][5] = 1;
assign rom[655][6] = 5;
assign rom[655][7] = 2;
assign rom[655][8] = -27;
assign rom[655][9] = 15;
assign rom[656][0] = -20;
assign rom[656][1] = 17;
assign rom[656][2] = -5;
assign rom[656][3] = -2;
assign rom[656][4] = -20;
assign rom[656][5] = 7;
assign rom[656][6] = -8;
assign rom[656][7] = 11;
assign rom[656][8] = -32;
assign rom[656][9] = 7;
assign rom[657][0] = -17;
assign rom[657][1] = 6;
assign rom[657][2] = -21;
assign rom[657][3] = 7;
assign rom[657][4] = -28;
assign rom[657][5] = 8;
assign rom[657][6] = -8;
assign rom[657][7] = 15;
assign rom[657][8] = -23;
assign rom[657][9] = 7;
assign rom[658][0] = -20;
assign rom[658][1] = 13;
assign rom[658][2] = -9;
assign rom[658][3] = -5;
assign rom[658][4] = -21;
assign rom[658][5] = 4;
assign rom[658][6] = -12;
assign rom[658][7] = 25;
assign rom[658][8] = -36;
assign rom[658][9] = 5;
assign rom[659][0] = -36;
assign rom[659][1] = -5;
assign rom[659][2] = -20;
assign rom[659][3] = 5;
assign rom[659][4] = -37;
assign rom[659][5] = 9;
assign rom[659][6] = 2;
assign rom[659][7] = 29;
assign rom[659][8] = -27;
assign rom[659][9] = 4;
assign rom[660][0] = -39;
assign rom[660][1] = -2;
assign rom[660][2] = -13;
assign rom[660][3] = 10;
assign rom[660][4] = -40;
assign rom[660][5] = 13;
assign rom[660][6] = -8;
assign rom[660][7] = 21;
assign rom[660][8] = -28;
assign rom[660][9] = 5;
assign rom[661][0] = -33;
assign rom[661][1] = 7;
assign rom[661][2] = -10;
assign rom[661][3] = 8;
assign rom[661][4] = -36;
assign rom[661][5] = 14;
assign rom[661][6] = -16;
assign rom[661][7] = 17;
assign rom[661][8] = -41;
assign rom[661][9] = 7;
assign rom[662][0] = -19;
assign rom[662][1] = 6;
assign rom[662][2] = -13;
assign rom[662][3] = 5;
assign rom[662][4] = -34;
assign rom[662][5] = -3;
assign rom[662][6] = -9;
assign rom[662][7] = 26;
assign rom[662][8] = -37;
assign rom[662][9] = 13;
assign rom[663][0] = -33;
assign rom[663][1] = -6;
assign rom[663][2] = -9;
assign rom[663][3] = 4;
assign rom[663][4] = -41;
assign rom[663][5] = 3;
assign rom[663][6] = -2;
assign rom[663][7] = 38;
assign rom[663][8] = -23;
assign rom[663][9] = 13;
assign rom[664][0] = -31;
assign rom[664][1] = 1;
assign rom[664][2] = -18;
assign rom[664][3] = -4;
assign rom[664][4] = -36;
assign rom[664][5] = -2;
assign rom[664][6] = -2;
assign rom[664][7] = 31;
assign rom[664][8] = -27;
assign rom[664][9] = 14;
assign rom[665][0] = -36;
assign rom[665][1] = 15;
assign rom[665][2] = -20;
assign rom[665][3] = -7;
assign rom[665][4] = -46;
assign rom[665][5] = 13;
assign rom[665][6] = -2;
assign rom[665][7] = 32;
assign rom[665][8] = -19;
assign rom[665][9] = 18;
assign rom[666][0] = -19;
assign rom[666][1] = 8;
assign rom[666][2] = -10;
assign rom[666][3] = -13;
assign rom[666][4] = -46;
assign rom[666][5] = 1;
assign rom[666][6] = -6;
assign rom[666][7] = 38;
assign rom[666][8] = -17;
assign rom[666][9] = 10;
assign rom[667][0] = -29;
assign rom[667][1] = 29;
assign rom[667][2] = -6;
assign rom[667][3] = -7;
assign rom[667][4] = -42;
assign rom[667][5] = -6;
assign rom[667][6] = 2;
assign rom[667][7] = 30;
assign rom[667][8] = -18;
assign rom[667][9] = 12;
assign rom[668][0] = -15;
assign rom[668][1] = 28;
assign rom[668][2] = -15;
assign rom[668][3] = -11;
assign rom[668][4] = -32;
assign rom[668][5] = 9;
assign rom[668][6] = -9;
assign rom[668][7] = 21;
assign rom[668][8] = -14;
assign rom[668][9] = 28;
assign rom[669][0] = -18;
assign rom[669][1] = 28;
assign rom[669][2] = -12;
assign rom[669][3] = -12;
assign rom[669][4] = -10;
assign rom[669][5] = 7;
assign rom[669][6] = 2;
assign rom[669][7] = 10;
assign rom[669][8] = -32;
assign rom[669][9] = 18;
assign rom[670][0] = -17;
assign rom[670][1] = 15;
assign rom[670][2] = -12;
assign rom[670][3] = -13;
assign rom[670][4] = -1;
assign rom[670][5] = 17;
assign rom[670][6] = 4;
assign rom[670][7] = 3;
assign rom[670][8] = -27;
assign rom[670][9] = 10;
assign rom[671][0] = -7;
assign rom[671][1] = 14;
assign rom[671][2] = 0;
assign rom[671][3] = -16;
assign rom[671][4] = 4;
assign rom[671][5] = 14;
assign rom[671][6] = -2;
assign rom[671][7] = 2;
assign rom[671][8] = -22;
assign rom[671][9] = 6;
assign rom[672][0] = -8;
assign rom[672][1] = 28;
assign rom[672][2] = -3;
assign rom[672][3] = -9;
assign rom[672][4] = 0;
assign rom[672][5] = 8;
assign rom[672][6] = -1;
assign rom[672][7] = 10;
assign rom[672][8] = -28;
assign rom[672][9] = 7;
assign rom[673][0] = 1;
assign rom[673][1] = 28;
assign rom[673][2] = -2;
assign rom[673][3] = -6;
assign rom[673][4] = 11;
assign rom[673][5] = 17;
assign rom[673][6] = 1;
assign rom[673][7] = 5;
assign rom[673][8] = -22;
assign rom[673][9] = 3;
assign rom[674][0] = -15;
assign rom[674][1] = 21;
assign rom[674][2] = -7;
assign rom[674][3] = -10;
assign rom[674][4] = 0;
assign rom[674][5] = 16;
assign rom[674][6] = 3;
assign rom[674][7] = 3;
assign rom[674][8] = -26;
assign rom[674][9] = 2;
assign rom[675][0] = -6;
assign rom[675][1] = 25;
assign rom[675][2] = -11;
assign rom[675][3] = -19;
assign rom[675][4] = 10;
assign rom[675][5] = 11;
assign rom[675][6] = -1;
assign rom[675][7] = 9;
assign rom[675][8] = -18;
assign rom[675][9] = 2;


endmodule

